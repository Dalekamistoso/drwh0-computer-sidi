library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4eac387",
    12 => x"86c0c64e",
    13 => x"49c4eac3",
    14 => x"48e0d0c3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e3e6",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"731e4f26",
    53 => x"029a721e",
    54 => x"c087e7c0",
    55 => x"724bc148",
    56 => x"87d106a9",
    57 => x"c9068272",
    58 => x"72837387",
    59 => x"87f401a9",
    60 => x"b2c187c3",
    61 => x"03a9723a",
    62 => x"07807389",
    63 => x"052b2ac1",
    64 => x"4b2687f3",
    65 => x"751e4f26",
    66 => x"714dc41e",
    67 => x"ff04a1b7",
    68 => x"c381c1b9",
    69 => x"b77207bd",
    70 => x"baff04a2",
    71 => x"bdc182c1",
    72 => x"87eefe07",
    73 => x"ff042dc1",
    74 => x"0780c1b8",
    75 => x"b9ff042d",
    76 => x"260781c1",
    77 => x"1e4f264d",
    78 => x"d4ff4811",
    79 => x"66c47808",
    80 => x"c888c148",
    81 => x"987058a6",
    82 => x"2687ed05",
    83 => x"d4ff1e4f",
    84 => x"78ffc348",
    85 => x"66c45168",
    86 => x"c888c148",
    87 => x"987058a6",
    88 => x"2687eb05",
    89 => x"1e731e4f",
    90 => x"c34bd4ff",
    91 => x"4a6b7bff",
    92 => x"6b7bffc3",
    93 => x"7232c849",
    94 => x"7bffc3b1",
    95 => x"31c84a6b",
    96 => x"ffc3b271",
    97 => x"c8496b7b",
    98 => x"71b17232",
    99 => x"2687c448",
   100 => x"264c264d",
   101 => x"0e4f264b",
   102 => x"5d5c5b5e",
   103 => x"ff4a710e",
   104 => x"49724cd4",
   105 => x"7199ffc3",
   106 => x"e0d0c37c",
   107 => x"87c805bf",
   108 => x"c94866d0",
   109 => x"58a6d430",
   110 => x"d84966d0",
   111 => x"99ffc329",
   112 => x"66d07c71",
   113 => x"c329d049",
   114 => x"7c7199ff",
   115 => x"c84966d0",
   116 => x"99ffc329",
   117 => x"66d07c71",
   118 => x"99ffc349",
   119 => x"49727c71",
   120 => x"ffc329d0",
   121 => x"6c7c7199",
   122 => x"fff0c94b",
   123 => x"abffc34d",
   124 => x"c387d005",
   125 => x"4b6c7cff",
   126 => x"c6028dc1",
   127 => x"abffc387",
   128 => x"7387f002",
   129 => x"87c7fe48",
   130 => x"ff49c01e",
   131 => x"ffc348d4",
   132 => x"c381c178",
   133 => x"04a9b7c8",
   134 => x"4f2687f1",
   135 => x"e71e731e",
   136 => x"dff8c487",
   137 => x"c01ec04b",
   138 => x"f7c1f0ff",
   139 => x"87e7fd49",
   140 => x"a8c186c4",
   141 => x"87eac005",
   142 => x"c348d4ff",
   143 => x"c0c178ff",
   144 => x"c0c0c0c0",
   145 => x"f0e1c01e",
   146 => x"fd49e9c1",
   147 => x"86c487c9",
   148 => x"ca059870",
   149 => x"48d4ff87",
   150 => x"c178ffc3",
   151 => x"fe87cb48",
   152 => x"8bc187e6",
   153 => x"87fdfe05",
   154 => x"e6fc48c0",
   155 => x"1e731e87",
   156 => x"c348d4ff",
   157 => x"4bd378ff",
   158 => x"ffc01ec0",
   159 => x"49c1c1f0",
   160 => x"c487d4fc",
   161 => x"05987086",
   162 => x"d4ff87ca",
   163 => x"78ffc348",
   164 => x"87cb48c1",
   165 => x"c187f1fd",
   166 => x"dbff058b",
   167 => x"fb48c087",
   168 => x"5e0e87f1",
   169 => x"ff0e5c5b",
   170 => x"dbfd4cd4",
   171 => x"1eeac687",
   172 => x"c1f0e1c0",
   173 => x"defb49c8",
   174 => x"c186c487",
   175 => x"87c802a8",
   176 => x"c087eafe",
   177 => x"87e2c148",
   178 => x"7087dafa",
   179 => x"ffffcf49",
   180 => x"a9eac699",
   181 => x"fe87c802",
   182 => x"48c087d3",
   183 => x"c387cbc1",
   184 => x"f1c07cff",
   185 => x"87f4fc4b",
   186 => x"c0029870",
   187 => x"1ec087eb",
   188 => x"c1f0ffc0",
   189 => x"defa49fa",
   190 => x"7086c487",
   191 => x"87d90598",
   192 => x"6c7cffc3",
   193 => x"7cffc349",
   194 => x"c17c7c7c",
   195 => x"c40299c0",
   196 => x"d548c187",
   197 => x"d148c087",
   198 => x"05abc287",
   199 => x"48c087c4",
   200 => x"8bc187c8",
   201 => x"87fdfe05",
   202 => x"e4f948c0",
   203 => x"1e731e87",
   204 => x"48e0d0c3",
   205 => x"4bc778c1",
   206 => x"c248d0ff",
   207 => x"87c8fb78",
   208 => x"c348d0ff",
   209 => x"c01ec078",
   210 => x"c0c1d0e5",
   211 => x"87c7f949",
   212 => x"a8c186c4",
   213 => x"4b87c105",
   214 => x"c505abc2",
   215 => x"c048c087",
   216 => x"8bc187f9",
   217 => x"87d0ff05",
   218 => x"c387f7fc",
   219 => x"7058e4d0",
   220 => x"87cd0598",
   221 => x"ffc01ec1",
   222 => x"49d0c1f0",
   223 => x"c487d8f8",
   224 => x"48d4ff86",
   225 => x"c478ffc3",
   226 => x"d0c387e0",
   227 => x"d0ff58e8",
   228 => x"ff78c248",
   229 => x"ffc348d4",
   230 => x"f748c178",
   231 => x"5e0e87f5",
   232 => x"0e5d5c5b",
   233 => x"ffc34a71",
   234 => x"4cd4ff4d",
   235 => x"d0ff7c75",
   236 => x"78c3c448",
   237 => x"1e727c75",
   238 => x"c1f0ffc0",
   239 => x"d6f749d8",
   240 => x"7086c487",
   241 => x"87c50298",
   242 => x"f0c048c0",
   243 => x"c37c7587",
   244 => x"c0c87cfe",
   245 => x"4966d41e",
   246 => x"c487dcf5",
   247 => x"757c7586",
   248 => x"d87c757c",
   249 => x"754be0da",
   250 => x"99496c7c",
   251 => x"c187c505",
   252 => x"87f3058b",
   253 => x"d0ff7c75",
   254 => x"c178c248",
   255 => x"87cff648",
   256 => x"4ad4ff1e",
   257 => x"c448d0ff",
   258 => x"ffc378d1",
   259 => x"0589c17a",
   260 => x"4f2687f8",
   261 => x"711e731e",
   262 => x"cdeec54b",
   263 => x"d4ff4adf",
   264 => x"78ffc348",
   265 => x"fec34868",
   266 => x"87c502a8",
   267 => x"ed058ac1",
   268 => x"059a7287",
   269 => x"48c087c5",
   270 => x"7387eac0",
   271 => x"87cc029b",
   272 => x"731e66c8",
   273 => x"87c5f449",
   274 => x"87c686c4",
   275 => x"fe4966c8",
   276 => x"d4ff87ee",
   277 => x"78ffc348",
   278 => x"059b7378",
   279 => x"d0ff87c5",
   280 => x"c178d048",
   281 => x"87ebf448",
   282 => x"711e731e",
   283 => x"ff4bc04a",
   284 => x"ffc348d4",
   285 => x"48d0ff78",
   286 => x"ff78c3c4",
   287 => x"ffc348d4",
   288 => x"c01e7278",
   289 => x"d1c1f0ff",
   290 => x"87cbf449",
   291 => x"987086c4",
   292 => x"c887cd05",
   293 => x"66cc1ec0",
   294 => x"87f8fd49",
   295 => x"4b7086c4",
   296 => x"c248d0ff",
   297 => x"f3487378",
   298 => x"5e0e87e9",
   299 => x"0e5d5c5b",
   300 => x"ffc01ec0",
   301 => x"49c9c1f0",
   302 => x"d287dcf3",
   303 => x"e8d0c31e",
   304 => x"87d0fd49",
   305 => x"4cc086c8",
   306 => x"b7d284c1",
   307 => x"87f804ac",
   308 => x"97e8d0c3",
   309 => x"c0c349bf",
   310 => x"a9c0c199",
   311 => x"87e7c005",
   312 => x"97efd0c3",
   313 => x"31d049bf",
   314 => x"97f0d0c3",
   315 => x"32c84abf",
   316 => x"d0c3b172",
   317 => x"4abf97f1",
   318 => x"cf4c71b1",
   319 => x"9cffffff",
   320 => x"34ca84c1",
   321 => x"c387e7c1",
   322 => x"bf97f1d0",
   323 => x"c631c149",
   324 => x"f2d0c399",
   325 => x"c74abf97",
   326 => x"b1722ab7",
   327 => x"97edd0c3",
   328 => x"cf4d4abf",
   329 => x"eed0c39d",
   330 => x"c34abf97",
   331 => x"c332ca9a",
   332 => x"bf97efd0",
   333 => x"7333c24b",
   334 => x"f0d0c3b2",
   335 => x"c34bbf97",
   336 => x"b7c69bc0",
   337 => x"c2b2732b",
   338 => x"7148c181",
   339 => x"c1497030",
   340 => x"70307548",
   341 => x"c14c724d",
   342 => x"c8947184",
   343 => x"06adb7c0",
   344 => x"34c187cc",
   345 => x"c0c82db7",
   346 => x"ff01adb7",
   347 => x"487487f4",
   348 => x"0e87dcf0",
   349 => x"5d5c5b5e",
   350 => x"c386f80e",
   351 => x"c048ced9",
   352 => x"c6d1c378",
   353 => x"fb49c01e",
   354 => x"86c487de",
   355 => x"c5059870",
   356 => x"c948c087",
   357 => x"4dc087ce",
   358 => x"fac07ec1",
   359 => x"c349bff2",
   360 => x"714afcd1",
   361 => x"c1eb4bc8",
   362 => x"05987087",
   363 => x"7ec087c2",
   364 => x"bfeefac0",
   365 => x"d8d2c349",
   366 => x"4bc8714a",
   367 => x"7087ebea",
   368 => x"87c20598",
   369 => x"026e7ec0",
   370 => x"c387fdc0",
   371 => x"4dbfccd8",
   372 => x"9fc4d9c3",
   373 => x"c5487ebf",
   374 => x"05a8ead6",
   375 => x"d8c387c7",
   376 => x"ce4dbfcc",
   377 => x"ca486e87",
   378 => x"02a8d5e9",
   379 => x"48c087c5",
   380 => x"c387f1c7",
   381 => x"751ec6d1",
   382 => x"87ecf949",
   383 => x"987086c4",
   384 => x"c087c505",
   385 => x"87dcc748",
   386 => x"bfeefac0",
   387 => x"d8d2c349",
   388 => x"4bc8714a",
   389 => x"7087d3e9",
   390 => x"87c80598",
   391 => x"48ced9c3",
   392 => x"87da78c1",
   393 => x"bff2fac0",
   394 => x"fcd1c349",
   395 => x"4bc8714a",
   396 => x"7087f7e8",
   397 => x"c5c00298",
   398 => x"c648c087",
   399 => x"d9c387e6",
   400 => x"49bf97c4",
   401 => x"05a9d5c1",
   402 => x"c387cdc0",
   403 => x"bf97c5d9",
   404 => x"a9eac249",
   405 => x"87c5c002",
   406 => x"c7c648c0",
   407 => x"c6d1c387",
   408 => x"487ebf97",
   409 => x"02a8e9c3",
   410 => x"6e87cec0",
   411 => x"a8ebc348",
   412 => x"87c5c002",
   413 => x"ebc548c0",
   414 => x"d1d1c387",
   415 => x"9949bf97",
   416 => x"87ccc005",
   417 => x"97d2d1c3",
   418 => x"a9c249bf",
   419 => x"87c5c002",
   420 => x"cfc548c0",
   421 => x"d3d1c387",
   422 => x"c348bf97",
   423 => x"7058cad9",
   424 => x"88c1484c",
   425 => x"58ced9c3",
   426 => x"97d4d1c3",
   427 => x"817549bf",
   428 => x"97d5d1c3",
   429 => x"32c84abf",
   430 => x"c37ea172",
   431 => x"6e48dbdd",
   432 => x"d6d1c378",
   433 => x"c848bf97",
   434 => x"d9c358a6",
   435 => x"c202bfce",
   436 => x"fac087d4",
   437 => x"c349bfee",
   438 => x"714ad8d2",
   439 => x"c9e64bc8",
   440 => x"02987087",
   441 => x"c087c5c0",
   442 => x"87f8c348",
   443 => x"bfc6d9c3",
   444 => x"efddc34c",
   445 => x"ebd1c35c",
   446 => x"c849bf97",
   447 => x"ead1c331",
   448 => x"a14abf97",
   449 => x"ecd1c349",
   450 => x"d04abf97",
   451 => x"49a17232",
   452 => x"97edd1c3",
   453 => x"32d84abf",
   454 => x"c449a172",
   455 => x"ddc39166",
   456 => x"c381bfdb",
   457 => x"c359e3dd",
   458 => x"bf97f3d1",
   459 => x"c332c84a",
   460 => x"bf97f2d1",
   461 => x"c34aa24b",
   462 => x"bf97f4d1",
   463 => x"7333d04b",
   464 => x"d1c34aa2",
   465 => x"4bbf97f5",
   466 => x"33d89bcf",
   467 => x"c34aa273",
   468 => x"c35ae7dd",
   469 => x"4abfe3dd",
   470 => x"92748ac2",
   471 => x"48e7ddc3",
   472 => x"c178a172",
   473 => x"d1c387ca",
   474 => x"49bf97d8",
   475 => x"d1c331c8",
   476 => x"4abf97d7",
   477 => x"d9c349a1",
   478 => x"d9c359d6",
   479 => x"c549bfd2",
   480 => x"81ffc731",
   481 => x"ddc329c9",
   482 => x"d1c359ef",
   483 => x"4abf97dd",
   484 => x"d1c332c8",
   485 => x"4bbf97dc",
   486 => x"66c44aa2",
   487 => x"c3826e92",
   488 => x"c35aebdd",
   489 => x"c048e3dd",
   490 => x"dfddc378",
   491 => x"78a17248",
   492 => x"48efddc3",
   493 => x"bfe3ddc3",
   494 => x"f3ddc378",
   495 => x"e7ddc348",
   496 => x"d9c378bf",
   497 => x"c002bfce",
   498 => x"487487c9",
   499 => x"7e7030c4",
   500 => x"c387c9c0",
   501 => x"48bfebdd",
   502 => x"7e7030c4",
   503 => x"48d2d9c3",
   504 => x"48c1786e",
   505 => x"4d268ef8",
   506 => x"4b264c26",
   507 => x"5e0e4f26",
   508 => x"0e5d5c5b",
   509 => x"d9c34a71",
   510 => x"cb02bfce",
   511 => x"c74b7287",
   512 => x"c14c722b",
   513 => x"87c99cff",
   514 => x"2bc84b72",
   515 => x"ffc34c72",
   516 => x"dbddc39c",
   517 => x"fac083bf",
   518 => x"02abbfea",
   519 => x"fac087d9",
   520 => x"d1c35bee",
   521 => x"49731ec6",
   522 => x"c487fdf0",
   523 => x"05987086",
   524 => x"48c087c5",
   525 => x"c387e6c0",
   526 => x"02bfced9",
   527 => x"497487d2",
   528 => x"d1c391c4",
   529 => x"4d6981c6",
   530 => x"ffffffcf",
   531 => x"87cb9dff",
   532 => x"91c24974",
   533 => x"81c6d1c3",
   534 => x"754d699f",
   535 => x"87c6fe48",
   536 => x"5c5b5e0e",
   537 => x"711e0e5d",
   538 => x"c11ec04d",
   539 => x"87e2d149",
   540 => x"4c7086c4",
   541 => x"c2c1029c",
   542 => x"d6d9c387",
   543 => x"ff49754a",
   544 => x"7087ccdf",
   545 => x"f2c00298",
   546 => x"754a7487",
   547 => x"ff4bcb49",
   548 => x"7087f1df",
   549 => x"e2c00298",
   550 => x"741ec087",
   551 => x"87c7029c",
   552 => x"c048a6c4",
   553 => x"c487c578",
   554 => x"78c148a6",
   555 => x"d04966c4",
   556 => x"86c487e0",
   557 => x"059c4c70",
   558 => x"7487fefe",
   559 => x"e5fc2648",
   560 => x"5b5e0e87",
   561 => x"f80e5d5c",
   562 => x"9b4b7186",
   563 => x"c087c505",
   564 => x"87d4c248",
   565 => x"c04da3c8",
   566 => x"0266d87d",
   567 => x"66d887c7",
   568 => x"c505bf97",
   569 => x"c148c087",
   570 => x"66d887fe",
   571 => x"87f0fd49",
   572 => x"026e7e70",
   573 => x"6e87efc1",
   574 => x"6981dc49",
   575 => x"da496e7d",
   576 => x"4ca3c481",
   577 => x"c37c699f",
   578 => x"02bfced9",
   579 => x"496e87d0",
   580 => x"699f81d4",
   581 => x"ffc04a49",
   582 => x"32d09aff",
   583 => x"4ac087c2",
   584 => x"6c484972",
   585 => x"c07c7080",
   586 => x"49a3cc7b",
   587 => x"a3d0796c",
   588 => x"c479c049",
   589 => x"78c048a6",
   590 => x"c44aa3d4",
   591 => x"91c84966",
   592 => x"c049a172",
   593 => x"c4796c41",
   594 => x"80c14866",
   595 => x"d058a6c8",
   596 => x"ff04a8b7",
   597 => x"4a6d87e2",
   598 => x"2ac72ac9",
   599 => x"49a3d4c2",
   600 => x"486e7972",
   601 => x"48c087c2",
   602 => x"f9f98ef8",
   603 => x"5b5e0e87",
   604 => x"710e5d5c",
   605 => x"eafac04c",
   606 => x"7478ff48",
   607 => x"cac1029c",
   608 => x"49a4c887",
   609 => x"c2c10269",
   610 => x"4a66d087",
   611 => x"d482496c",
   612 => x"66d05aa6",
   613 => x"d9c3b94d",
   614 => x"ff4abfca",
   615 => x"719972ba",
   616 => x"e4c00299",
   617 => x"4ba4c487",
   618 => x"c1f9496b",
   619 => x"c37b7087",
   620 => x"49bfc6d9",
   621 => x"7c71816c",
   622 => x"d9c3b975",
   623 => x"ff4abfca",
   624 => x"719972ba",
   625 => x"dcff0599",
   626 => x"f87c7587",
   627 => x"731e87d8",
   628 => x"9b4b711e",
   629 => x"c887c702",
   630 => x"056949a3",
   631 => x"48c087c5",
   632 => x"c387ebc0",
   633 => x"4abfdfdd",
   634 => x"6949a3c4",
   635 => x"c389c249",
   636 => x"91bfc6d9",
   637 => x"c34aa271",
   638 => x"49bfcad9",
   639 => x"a271996b",
   640 => x"1e66c84a",
   641 => x"dfe94972",
   642 => x"7086c487",
   643 => x"d9f74849",
   644 => x"1e731e87",
   645 => x"029b4b71",
   646 => x"a3c887c7",
   647 => x"c5056949",
   648 => x"c048c087",
   649 => x"ddc387eb",
   650 => x"c44abfdf",
   651 => x"496949a3",
   652 => x"d9c389c2",
   653 => x"7191bfc6",
   654 => x"d9c34aa2",
   655 => x"6b49bfca",
   656 => x"4aa27199",
   657 => x"721e66c8",
   658 => x"87d2e549",
   659 => x"497086c4",
   660 => x"87d6f648",
   661 => x"5c5b5e0e",
   662 => x"86f80e5d",
   663 => x"a6c44b71",
   664 => x"c878ff48",
   665 => x"4d6949a3",
   666 => x"a3d44cc0",
   667 => x"c849744a",
   668 => x"49a17291",
   669 => x"66d84969",
   670 => x"70887148",
   671 => x"a966d87e",
   672 => x"6e87ca01",
   673 => x"87c506ad",
   674 => x"6e5ca6c8",
   675 => x"d084c14d",
   676 => x"ff04acb7",
   677 => x"66c487d4",
   678 => x"f58ef848",
   679 => x"5e0e87c8",
   680 => x"0e5d5c5b",
   681 => x"a6c886ec",
   682 => x"48a6c859",
   683 => x"ffffffc1",
   684 => x"c478ffff",
   685 => x"c078ff80",
   686 => x"c44cc04d",
   687 => x"83d44b66",
   688 => x"91c84974",
   689 => x"7549a173",
   690 => x"7392c84a",
   691 => x"49697ea2",
   692 => x"d489bf6e",
   693 => x"ad7459a6",
   694 => x"d087c605",
   695 => x"bf6e48a6",
   696 => x"4866d078",
   697 => x"04a8b7c0",
   698 => x"66d087cf",
   699 => x"a966c849",
   700 => x"d087c603",
   701 => x"a6cc5ca6",
   702 => x"d084c159",
   703 => x"fe04acb7",
   704 => x"85c187f9",
   705 => x"04adb7d0",
   706 => x"cc87eefe",
   707 => x"8eec4866",
   708 => x"0e87d3f3",
   709 => x"0e5c5b5e",
   710 => x"4cc04b71",
   711 => x"6949a3c8",
   712 => x"7429c449",
   713 => x"1e71914a",
   714 => x"87d44973",
   715 => x"84c186c4",
   716 => x"04acb7d0",
   717 => x"1ec087e6",
   718 => x"87c44973",
   719 => x"87e8f226",
   720 => x"5c5b5e0e",
   721 => x"86f00e5d",
   722 => x"e0c04b71",
   723 => x"2cc94c66",
   724 => x"c3029b73",
   725 => x"a3c887e1",
   726 => x"c3026949",
   727 => x"a3d087d9",
   728 => x"66e0c049",
   729 => x"ac7e6b79",
   730 => x"87cbc302",
   731 => x"bfcad9c3",
   732 => x"71b9ff49",
   733 => x"719a744a",
   734 => x"cc986e48",
   735 => x"a3c458a6",
   736 => x"48a6c44d",
   737 => x"66c8786d",
   738 => x"87c505aa",
   739 => x"d1c27b74",
   740 => x"731e7287",
   741 => x"87fcfa49",
   742 => x"7e7086c4",
   743 => x"a8b7c048",
   744 => x"d487d004",
   745 => x"496e4aa3",
   746 => x"a17291c8",
   747 => x"697b2149",
   748 => x"c087c77d",
   749 => x"49a3cc7b",
   750 => x"66c87d69",
   751 => x"fa49731e",
   752 => x"86c487d2",
   753 => x"d4c27e70",
   754 => x"a6cc49a3",
   755 => x"c8786948",
   756 => x"66cc4866",
   757 => x"87c906a8",
   758 => x"b7c0486e",
   759 => x"e0c004a8",
   760 => x"c0486e87",
   761 => x"c004a8b7",
   762 => x"a3d487ec",
   763 => x"c8496e4a",
   764 => x"49a17291",
   765 => x"694866c8",
   766 => x"cc497088",
   767 => x"d506a966",
   768 => x"fa497387",
   769 => x"497087d8",
   770 => x"c84aa3d4",
   771 => x"49a17291",
   772 => x"c44166c8",
   773 => x"8c6b7966",
   774 => x"731e4974",
   775 => x"87cdf549",
   776 => x"e0c086c4",
   777 => x"ffc74966",
   778 => x"87cb0299",
   779 => x"1ec6d1c3",
   780 => x"d9f64973",
   781 => x"f086c487",
   782 => x"87eaee8e",
   783 => x"711e731e",
   784 => x"c0029b4b",
   785 => x"ddc387e4",
   786 => x"4a735bf3",
   787 => x"d9c38ac2",
   788 => x"9249bfc6",
   789 => x"bfdfddc3",
   790 => x"c3807248",
   791 => x"7158f7dd",
   792 => x"c330c448",
   793 => x"c058d6d9",
   794 => x"ddc387ed",
   795 => x"ddc348ef",
   796 => x"c378bfe3",
   797 => x"c348f3dd",
   798 => x"78bfe7dd",
   799 => x"bfced9c3",
   800 => x"c387c902",
   801 => x"49bfc6d9",
   802 => x"87c731c4",
   803 => x"bfebddc3",
   804 => x"c331c449",
   805 => x"ed59d6d9",
   806 => x"5e0e87d0",
   807 => x"710e5c5b",
   808 => x"724bc04a",
   809 => x"e1c0029a",
   810 => x"49a2da87",
   811 => x"c34b699f",
   812 => x"02bfced9",
   813 => x"a2d487cf",
   814 => x"49699f49",
   815 => x"ffffc04c",
   816 => x"c234d09c",
   817 => x"744cc087",
   818 => x"4973b349",
   819 => x"ec87edfd",
   820 => x"5e0e87d6",
   821 => x"0e5d5c5b",
   822 => x"4a7186f4",
   823 => x"9a727ec0",
   824 => x"c387d802",
   825 => x"c048c2d1",
   826 => x"fad0c378",
   827 => x"f3ddc348",
   828 => x"d0c378bf",
   829 => x"ddc348fe",
   830 => x"c378bfef",
   831 => x"c048e3d9",
   832 => x"d2d9c350",
   833 => x"d1c349bf",
   834 => x"714abfc2",
   835 => x"c0c403aa",
   836 => x"cf497287",
   837 => x"e1c00599",
   838 => x"c6d1c387",
   839 => x"fad0c31e",
   840 => x"d0c349bf",
   841 => x"a1c148fa",
   842 => x"dcff7178",
   843 => x"86c487fa",
   844 => x"48e6fac0",
   845 => x"78c6d1c3",
   846 => x"fac087cc",
   847 => x"c048bfe6",
   848 => x"fac080e0",
   849 => x"d1c358ea",
   850 => x"c148bfc2",
   851 => x"c6d1c380",
   852 => x"0ea62758",
   853 => x"97bf0000",
   854 => x"029d4dbf",
   855 => x"c387e2c2",
   856 => x"c202ade5",
   857 => x"fac087db",
   858 => x"cb4bbfe6",
   859 => x"4c1149a3",
   860 => x"c105accf",
   861 => x"497587d2",
   862 => x"89c199df",
   863 => x"d9c391cd",
   864 => x"a3c181d6",
   865 => x"c351124a",
   866 => x"51124aa3",
   867 => x"124aa3c5",
   868 => x"4aa3c751",
   869 => x"a3c95112",
   870 => x"ce51124a",
   871 => x"51124aa3",
   872 => x"124aa3d0",
   873 => x"4aa3d251",
   874 => x"a3d45112",
   875 => x"d651124a",
   876 => x"51124aa3",
   877 => x"124aa3d8",
   878 => x"4aa3dc51",
   879 => x"a3de5112",
   880 => x"c151124a",
   881 => x"87f9c07e",
   882 => x"99c84974",
   883 => x"87eac005",
   884 => x"99d04974",
   885 => x"dc87d005",
   886 => x"cac00266",
   887 => x"dc497387",
   888 => x"98700f66",
   889 => x"6e87d302",
   890 => x"87c6c005",
   891 => x"48d6d9c3",
   892 => x"fac050c0",
   893 => x"c248bfe6",
   894 => x"d9c387e7",
   895 => x"50c048e3",
   896 => x"d2d9c37e",
   897 => x"d1c349bf",
   898 => x"714abfc2",
   899 => x"c0fc04aa",
   900 => x"f3ddc387",
   901 => x"c8c005bf",
   902 => x"ced9c387",
   903 => x"fec102bf",
   904 => x"eafac087",
   905 => x"c378ff48",
   906 => x"49bffed0",
   907 => x"7087ffe6",
   908 => x"c2d1c349",
   909 => x"48a6c459",
   910 => x"bffed0c3",
   911 => x"ced9c378",
   912 => x"d8c002bf",
   913 => x"4966c487",
   914 => x"ffffffcf",
   915 => x"02a999f8",
   916 => x"c087c5c0",
   917 => x"87e1c04d",
   918 => x"dcc04dc1",
   919 => x"4966c487",
   920 => x"99f8ffcf",
   921 => x"c8c002a9",
   922 => x"48a6c887",
   923 => x"c5c078c0",
   924 => x"48a6c887",
   925 => x"66c878c1",
   926 => x"059d754d",
   927 => x"c487e0c0",
   928 => x"89c24966",
   929 => x"bfc6d9c3",
   930 => x"ddc3914a",
   931 => x"c34abfdf",
   932 => x"7248fad0",
   933 => x"d1c378a1",
   934 => x"78c048c2",
   935 => x"c087e2f9",
   936 => x"e58ef448",
   937 => x"000087c0",
   938 => x"ffff0000",
   939 => x"0eb6ffff",
   940 => x"0ebf0000",
   941 => x"41460000",
   942 => x"20323354",
   943 => x"46002020",
   944 => x"36315441",
   945 => x"00202020",
   946 => x"48d4ff1e",
   947 => x"6878ffc3",
   948 => x"1e4f2648",
   949 => x"c348d4ff",
   950 => x"d0ff78ff",
   951 => x"78e1c848",
   952 => x"d448d4ff",
   953 => x"f7ddc378",
   954 => x"bfd4ff48",
   955 => x"1e4f2650",
   956 => x"c048d0ff",
   957 => x"4f2678e0",
   958 => x"87ccff1e",
   959 => x"02994970",
   960 => x"fbc087c6",
   961 => x"87f105a9",
   962 => x"4f264871",
   963 => x"5c5b5e0e",
   964 => x"c04b710e",
   965 => x"87f0fe4c",
   966 => x"02994970",
   967 => x"c087f9c0",
   968 => x"c002a9ec",
   969 => x"fbc087f2",
   970 => x"ebc002a9",
   971 => x"b766cc87",
   972 => x"87c703ac",
   973 => x"c20266d0",
   974 => x"71537187",
   975 => x"87c20299",
   976 => x"c3fe84c1",
   977 => x"99497087",
   978 => x"c087cd02",
   979 => x"c702a9ec",
   980 => x"a9fbc087",
   981 => x"87d5ff05",
   982 => x"c30266d0",
   983 => x"7b97c087",
   984 => x"05a9ecc0",
   985 => x"4a7487c4",
   986 => x"4a7487c5",
   987 => x"728a0ac0",
   988 => x"2687c248",
   989 => x"264c264d",
   990 => x"1e4f264b",
   991 => x"7087c9fd",
   992 => x"b7f0c049",
   993 => x"87ca04a9",
   994 => x"a9b7f9c0",
   995 => x"c087c301",
   996 => x"c1c189f0",
   997 => x"ca04a9b7",
   998 => x"b7dac187",
   999 => x"87c301a9",
  1000 => x"c189f7c0",
  1001 => x"04a9b7e1",
  1002 => x"fac187ca",
  1003 => x"c301a9b7",
  1004 => x"89fdc087",
  1005 => x"4f264871",
  1006 => x"5c5b5e0e",
  1007 => x"ff4a710e",
  1008 => x"49724cd4",
  1009 => x"7087eac0",
  1010 => x"c2029b4b",
  1011 => x"ff8bc187",
  1012 => x"c5c848d0",
  1013 => x"7cd5c178",
  1014 => x"31c64973",
  1015 => x"97d5ccc3",
  1016 => x"71484abf",
  1017 => x"ff7c70b0",
  1018 => x"78c448d0",
  1019 => x"c4fe4873",
  1020 => x"5b5e0e87",
  1021 => x"f80e5d5c",
  1022 => x"c04c7186",
  1023 => x"87d3fb7e",
  1024 => x"c2c14bc0",
  1025 => x"49bf97de",
  1026 => x"cf04a9c0",
  1027 => x"87e8fb87",
  1028 => x"c2c183c1",
  1029 => x"49bf97de",
  1030 => x"87f106ab",
  1031 => x"97dec2c1",
  1032 => x"87cf02bf",
  1033 => x"7087e1fa",
  1034 => x"c6029949",
  1035 => x"a9ecc087",
  1036 => x"c087f105",
  1037 => x"87d0fa4b",
  1038 => x"cbfa4d70",
  1039 => x"58a6c887",
  1040 => x"7087c5fa",
  1041 => x"c883c14a",
  1042 => x"699749a4",
  1043 => x"c702ad49",
  1044 => x"adffc087",
  1045 => x"87e7c005",
  1046 => x"9749a4c9",
  1047 => x"66c44969",
  1048 => x"87c702a9",
  1049 => x"a8ffc048",
  1050 => x"ca87d405",
  1051 => x"699749a4",
  1052 => x"c602aa49",
  1053 => x"aaffc087",
  1054 => x"c187c405",
  1055 => x"c087d07e",
  1056 => x"c602adec",
  1057 => x"adfbc087",
  1058 => x"c087c405",
  1059 => x"6e7ec14b",
  1060 => x"87e1fe02",
  1061 => x"7387d8f9",
  1062 => x"fb8ef848",
  1063 => x"0e0087d5",
  1064 => x"5d5c5b5e",
  1065 => x"4b711e0e",
  1066 => x"ab4d4cc0",
  1067 => x"87e8c004",
  1068 => x"1ef1ffc0",
  1069 => x"c4029d75",
  1070 => x"c24ac087",
  1071 => x"724ac187",
  1072 => x"87cef049",
  1073 => x"7e7086c4",
  1074 => x"056e84c1",
  1075 => x"4c7387c2",
  1076 => x"ac7385c1",
  1077 => x"87d8ff06",
  1078 => x"2626486e",
  1079 => x"264c264d",
  1080 => x"0e4f264b",
  1081 => x"5d5c5b5e",
  1082 => x"4c711e0e",
  1083 => x"c391de49",
  1084 => x"714dd1de",
  1085 => x"026d9785",
  1086 => x"c387ddc1",
  1087 => x"4abffcdd",
  1088 => x"49728274",
  1089 => x"7087d8fe",
  1090 => x"c0026e7e",
  1091 => x"dec387f3",
  1092 => x"4a6e4bc4",
  1093 => x"fefe49cb",
  1094 => x"4b7487ce",
  1095 => x"e8c193cb",
  1096 => x"83c483d3",
  1097 => x"7bdcc5c1",
  1098 => x"c8c14974",
  1099 => x"7b7587f2",
  1100 => x"97d0dec3",
  1101 => x"c31e49bf",
  1102 => x"c249c4de",
  1103 => x"c487dfc6",
  1104 => x"c1497486",
  1105 => x"c087d9c8",
  1106 => x"f8c9c149",
  1107 => x"f8ddc387",
  1108 => x"c178c048",
  1109 => x"87cfdd49",
  1110 => x"87fffd26",
  1111 => x"64616f4c",
  1112 => x"2e676e69",
  1113 => x"0e002e2e",
  1114 => x"0e5c5b5e",
  1115 => x"c34a4b71",
  1116 => x"82bffcdd",
  1117 => x"e6fc4972",
  1118 => x"9c4c7087",
  1119 => x"4987c402",
  1120 => x"c387d7ec",
  1121 => x"c048fcdd",
  1122 => x"dc49c178",
  1123 => x"ccfd87d9",
  1124 => x"5b5e0e87",
  1125 => x"f40e5d5c",
  1126 => x"c6d1c386",
  1127 => x"c44cc04d",
  1128 => x"78c048a6",
  1129 => x"bffcddc3",
  1130 => x"06a9c049",
  1131 => x"c387c1c1",
  1132 => x"9848c6d1",
  1133 => x"87f8c002",
  1134 => x"1ef1ffc0",
  1135 => x"c70266c8",
  1136 => x"48a6c487",
  1137 => x"87c578c0",
  1138 => x"c148a6c4",
  1139 => x"4966c478",
  1140 => x"c487ffeb",
  1141 => x"c14d7086",
  1142 => x"4866c484",
  1143 => x"a6c880c1",
  1144 => x"fcddc358",
  1145 => x"03ac49bf",
  1146 => x"9d7587c6",
  1147 => x"87c8ff05",
  1148 => x"9d754cc0",
  1149 => x"87e0c302",
  1150 => x"1ef1ffc0",
  1151 => x"c70266c8",
  1152 => x"48a6cc87",
  1153 => x"87c578c0",
  1154 => x"c148a6cc",
  1155 => x"4966cc78",
  1156 => x"c487ffea",
  1157 => x"6e7e7086",
  1158 => x"87e9c202",
  1159 => x"81cb496e",
  1160 => x"d0496997",
  1161 => x"d6c10299",
  1162 => x"e7c5c187",
  1163 => x"cb49744a",
  1164 => x"d3e8c191",
  1165 => x"c8797281",
  1166 => x"51ffc381",
  1167 => x"91de4974",
  1168 => x"4dd1dec3",
  1169 => x"c1c28571",
  1170 => x"a5c17d97",
  1171 => x"51e0c049",
  1172 => x"97d6d9c3",
  1173 => x"87d202bf",
  1174 => x"a5c284c1",
  1175 => x"d6d9c34b",
  1176 => x"fe49db4a",
  1177 => x"c187c1f9",
  1178 => x"a5cd87db",
  1179 => x"c151c049",
  1180 => x"4ba5c284",
  1181 => x"49cb4a6e",
  1182 => x"87ecf8fe",
  1183 => x"c187c6c1",
  1184 => x"744ae3c3",
  1185 => x"c191cb49",
  1186 => x"7281d3e8",
  1187 => x"d6d9c379",
  1188 => x"d802bf97",
  1189 => x"de497487",
  1190 => x"c384c191",
  1191 => x"714bd1de",
  1192 => x"d6d9c383",
  1193 => x"fe49dd4a",
  1194 => x"d887fdf7",
  1195 => x"de4b7487",
  1196 => x"d1dec393",
  1197 => x"49a3cb83",
  1198 => x"84c151c0",
  1199 => x"cb4a6e73",
  1200 => x"e3f7fe49",
  1201 => x"4866c487",
  1202 => x"a6c880c1",
  1203 => x"03acc758",
  1204 => x"6e87c5c0",
  1205 => x"87e0fc05",
  1206 => x"8ef44874",
  1207 => x"1e87fcf7",
  1208 => x"4b711e73",
  1209 => x"c191cb49",
  1210 => x"c881d3e8",
  1211 => x"ccc34aa1",
  1212 => x"501248d5",
  1213 => x"c14aa1c9",
  1214 => x"1248dec2",
  1215 => x"c381ca50",
  1216 => x"1148d0de",
  1217 => x"d0dec350",
  1218 => x"1e49bf97",
  1219 => x"ffc149c0",
  1220 => x"ddc387cc",
  1221 => x"78de48f8",
  1222 => x"cad649c1",
  1223 => x"fef62687",
  1224 => x"4a711e87",
  1225 => x"c191cb49",
  1226 => x"c881d3e8",
  1227 => x"c3481181",
  1228 => x"c358fcdd",
  1229 => x"c048fcdd",
  1230 => x"d549c178",
  1231 => x"4f2687e9",
  1232 => x"c149c01e",
  1233 => x"2687fec1",
  1234 => x"99711e4f",
  1235 => x"c187d202",
  1236 => x"c048e8e9",
  1237 => x"c180f750",
  1238 => x"c140e1cc",
  1239 => x"ce78cce8",
  1240 => x"e4e9c187",
  1241 => x"c5e8c148",
  1242 => x"c180fc78",
  1243 => x"2678c0cd",
  1244 => x"5b5e0e4f",
  1245 => x"4c710e5c",
  1246 => x"c192cb4a",
  1247 => x"c882d3e8",
  1248 => x"a2c949a2",
  1249 => x"4b6b974b",
  1250 => x"4969971e",
  1251 => x"1282ca1e",
  1252 => x"f7eac049",
  1253 => x"d449c087",
  1254 => x"497487cd",
  1255 => x"87c0ffc0",
  1256 => x"f8f48ef8",
  1257 => x"1e731e87",
  1258 => x"ff494b71",
  1259 => x"497387c3",
  1260 => x"c087fefe",
  1261 => x"ccc0c149",
  1262 => x"87e3f487",
  1263 => x"711e731e",
  1264 => x"4aa3c64b",
  1265 => x"c187db02",
  1266 => x"87d6028a",
  1267 => x"dac1028a",
  1268 => x"c0028a87",
  1269 => x"028a87fc",
  1270 => x"8a87e1c0",
  1271 => x"c187cb02",
  1272 => x"49c787db",
  1273 => x"c187fafc",
  1274 => x"ddc387de",
  1275 => x"c102bffc",
  1276 => x"c14887cb",
  1277 => x"c0dec388",
  1278 => x"87c1c158",
  1279 => x"bfc0dec3",
  1280 => x"87f9c002",
  1281 => x"bffcddc3",
  1282 => x"c380c148",
  1283 => x"c058c0de",
  1284 => x"ddc387eb",
  1285 => x"c649bffc",
  1286 => x"c0dec389",
  1287 => x"a9b7c059",
  1288 => x"c387da03",
  1289 => x"c048fcdd",
  1290 => x"c387d278",
  1291 => x"02bfc0de",
  1292 => x"ddc387cb",
  1293 => x"c648bffc",
  1294 => x"c0dec380",
  1295 => x"d149c058",
  1296 => x"497387e5",
  1297 => x"87d8fcc0",
  1298 => x"0e87d4f2",
  1299 => x"0e5c5b5e",
  1300 => x"66cc4c71",
  1301 => x"cb4b741e",
  1302 => x"d3e8c193",
  1303 => x"4aa3c483",
  1304 => x"f1fe496a",
  1305 => x"cbc187d2",
  1306 => x"a3c87bdf",
  1307 => x"5166d449",
  1308 => x"d849a3c9",
  1309 => x"a3ca5166",
  1310 => x"5166dc49",
  1311 => x"87ddf126",
  1312 => x"5c5b5e0e",
  1313 => x"d0ff0e5d",
  1314 => x"59a6d886",
  1315 => x"c048a6c4",
  1316 => x"c180c478",
  1317 => x"c47866c4",
  1318 => x"c478c180",
  1319 => x"c378c180",
  1320 => x"c148c0de",
  1321 => x"f8ddc378",
  1322 => x"a8de48bf",
  1323 => x"f387cb05",
  1324 => x"497087df",
  1325 => x"ce59a6c8",
  1326 => x"d6e887f6",
  1327 => x"87f8e887",
  1328 => x"7087c5e8",
  1329 => x"acfbc04c",
  1330 => x"87d0c102",
  1331 => x"c10566d4",
  1332 => x"1ec087c2",
  1333 => x"c11ec11e",
  1334 => x"c01ef6e9",
  1335 => x"87ebfd49",
  1336 => x"4a66d0c1",
  1337 => x"496a82c4",
  1338 => x"517481c7",
  1339 => x"1ed81ec1",
  1340 => x"81c8496a",
  1341 => x"d887d5e8",
  1342 => x"66c4c186",
  1343 => x"01a8c048",
  1344 => x"a6c487c7",
  1345 => x"ce78c148",
  1346 => x"66c4c187",
  1347 => x"cc88c148",
  1348 => x"87c358a6",
  1349 => x"cc87e1e7",
  1350 => x"78c248a6",
  1351 => x"cd029c74",
  1352 => x"66c487ca",
  1353 => x"66c8c148",
  1354 => x"ffcc03a8",
  1355 => x"48a6d887",
  1356 => x"d3e678c0",
  1357 => x"c14c7087",
  1358 => x"c205acd0",
  1359 => x"66d887d6",
  1360 => x"87f7e87e",
  1361 => x"a6dc4970",
  1362 => x"87fce559",
  1363 => x"ecc04c70",
  1364 => x"eac105ac",
  1365 => x"4966c487",
  1366 => x"c0c191cb",
  1367 => x"a1c48166",
  1368 => x"c84d6a4a",
  1369 => x"66d84aa1",
  1370 => x"e1ccc152",
  1371 => x"87d8e579",
  1372 => x"029c4c70",
  1373 => x"fbc087d8",
  1374 => x"87d202ac",
  1375 => x"c7e55574",
  1376 => x"9c4c7087",
  1377 => x"c087c702",
  1378 => x"ff05acfb",
  1379 => x"e0c087ee",
  1380 => x"55c1c255",
  1381 => x"d47d97c0",
  1382 => x"a96e4966",
  1383 => x"c487db05",
  1384 => x"66c84866",
  1385 => x"87ca04a8",
  1386 => x"c14866c4",
  1387 => x"58a6c880",
  1388 => x"66c887c8",
  1389 => x"cc88c148",
  1390 => x"cbe458a6",
  1391 => x"c14c7087",
  1392 => x"c805acd0",
  1393 => x"4866d087",
  1394 => x"a6d480c1",
  1395 => x"acd0c158",
  1396 => x"87eafd02",
  1397 => x"d448a6dc",
  1398 => x"66d87866",
  1399 => x"a866dc48",
  1400 => x"87dac905",
  1401 => x"48a6e0c0",
  1402 => x"c478f0c0",
  1403 => x"7866cc80",
  1404 => x"78c080c4",
  1405 => x"c048747e",
  1406 => x"f0c088fb",
  1407 => x"987058a6",
  1408 => x"87d5c802",
  1409 => x"c088cb48",
  1410 => x"7058a6f0",
  1411 => x"e9c00298",
  1412 => x"88c94887",
  1413 => x"58a6f0c0",
  1414 => x"c3029870",
  1415 => x"c44887e1",
  1416 => x"a6f0c088",
  1417 => x"02987058",
  1418 => x"c14887d6",
  1419 => x"a6f0c088",
  1420 => x"02987058",
  1421 => x"c787c8c3",
  1422 => x"e0c087d9",
  1423 => x"78c048a6",
  1424 => x"c14866cc",
  1425 => x"58a6d080",
  1426 => x"7087fde1",
  1427 => x"acecc04c",
  1428 => x"c087d502",
  1429 => x"c60266e0",
  1430 => x"a6e4c087",
  1431 => x"7487c95c",
  1432 => x"88f0c048",
  1433 => x"58a6e8c0",
  1434 => x"02acecc0",
  1435 => x"d7e187cc",
  1436 => x"c04c7087",
  1437 => x"ff05acec",
  1438 => x"e0c087f4",
  1439 => x"66d41e66",
  1440 => x"ecc01e49",
  1441 => x"e9c11e66",
  1442 => x"66d41ef6",
  1443 => x"87fbf649",
  1444 => x"1eca1ec0",
  1445 => x"cb4966dc",
  1446 => x"66d8c191",
  1447 => x"48a6d881",
  1448 => x"d878a1c4",
  1449 => x"e149bf66",
  1450 => x"86d887e2",
  1451 => x"06a8b7c0",
  1452 => x"c187c7c1",
  1453 => x"c81ede1e",
  1454 => x"e149bf66",
  1455 => x"86c887ce",
  1456 => x"c0484970",
  1457 => x"e4c08808",
  1458 => x"b7c058a6",
  1459 => x"e9c006a8",
  1460 => x"66e0c087",
  1461 => x"a8b7dd48",
  1462 => x"6e87df03",
  1463 => x"e0c049bf",
  1464 => x"e0c08166",
  1465 => x"c1496651",
  1466 => x"81bf6e81",
  1467 => x"c051c1c2",
  1468 => x"c24966e0",
  1469 => x"81bf6e81",
  1470 => x"7ec151c0",
  1471 => x"e187dac4",
  1472 => x"e4c087f9",
  1473 => x"f2e158a6",
  1474 => x"a6e8c087",
  1475 => x"a8ecc058",
  1476 => x"87cbc005",
  1477 => x"48a6e4c0",
  1478 => x"7866e0c0",
  1479 => x"ff87c4c0",
  1480 => x"c487e5de",
  1481 => x"91cb4966",
  1482 => x"4866c0c1",
  1483 => x"7e708071",
  1484 => x"81c8496e",
  1485 => x"82ca4a6e",
  1486 => x"5266e0c0",
  1487 => x"4a66e4c0",
  1488 => x"e0c082c1",
  1489 => x"48c18a66",
  1490 => x"4a703072",
  1491 => x"97728ac1",
  1492 => x"49699779",
  1493 => x"66e4c01e",
  1494 => x"87f2da49",
  1495 => x"f0c086c4",
  1496 => x"496e58a6",
  1497 => x"4d6981c4",
  1498 => x"d84866dc",
  1499 => x"c002a866",
  1500 => x"a6d887c8",
  1501 => x"c078c048",
  1502 => x"a6d887c5",
  1503 => x"d878c148",
  1504 => x"e0c01e66",
  1505 => x"ff49751e",
  1506 => x"c887c1de",
  1507 => x"c04c7086",
  1508 => x"c106acb7",
  1509 => x"857487d4",
  1510 => x"7449e0c0",
  1511 => x"c14b7589",
  1512 => x"714ae4e2",
  1513 => x"87c0e4fe",
  1514 => x"e8c085c2",
  1515 => x"80c14866",
  1516 => x"58a6ecc0",
  1517 => x"4966ecc0",
  1518 => x"a97081c1",
  1519 => x"87c8c002",
  1520 => x"c048a6d8",
  1521 => x"87c5c078",
  1522 => x"c148a6d8",
  1523 => x"1e66d878",
  1524 => x"c049a4c2",
  1525 => x"887148e0",
  1526 => x"751e4970",
  1527 => x"ebdcff49",
  1528 => x"c086c887",
  1529 => x"ff01a8b7",
  1530 => x"e8c087c0",
  1531 => x"d1c00266",
  1532 => x"c9496e87",
  1533 => x"66e8c081",
  1534 => x"c1486e51",
  1535 => x"c078f1cd",
  1536 => x"496e87cc",
  1537 => x"51c281c9",
  1538 => x"cec1486e",
  1539 => x"7ec178e5",
  1540 => x"ff87c6c0",
  1541 => x"7087e1db",
  1542 => x"c0026e4c",
  1543 => x"66c487f5",
  1544 => x"a866c848",
  1545 => x"87cbc004",
  1546 => x"c14866c4",
  1547 => x"58a6c880",
  1548 => x"c887e0c0",
  1549 => x"88c14866",
  1550 => x"c058a6cc",
  1551 => x"c6c187d5",
  1552 => x"c8c005ac",
  1553 => x"4866cc87",
  1554 => x"a6d080c1",
  1555 => x"e7daff58",
  1556 => x"d04c7087",
  1557 => x"80c14866",
  1558 => x"7458a6d4",
  1559 => x"cbc0029c",
  1560 => x"4866c487",
  1561 => x"a866c8c1",
  1562 => x"87c1f304",
  1563 => x"87ffd9ff",
  1564 => x"c74866c4",
  1565 => x"e5c003a8",
  1566 => x"c0dec387",
  1567 => x"c478c048",
  1568 => x"91cb4966",
  1569 => x"8166c0c1",
  1570 => x"6a4aa1c4",
  1571 => x"7952c04a",
  1572 => x"c14866c4",
  1573 => x"58a6c880",
  1574 => x"ff04a8c7",
  1575 => x"d0ff87db",
  1576 => x"87f7e08e",
  1577 => x"1e00203a",
  1578 => x"4b711e73",
  1579 => x"87c6029b",
  1580 => x"48fcddc3",
  1581 => x"1ec778c0",
  1582 => x"bffcddc3",
  1583 => x"e8c11e49",
  1584 => x"ddc31ed3",
  1585 => x"ee49bff8",
  1586 => x"86cc87f6",
  1587 => x"bff8ddc3",
  1588 => x"87f5e949",
  1589 => x"c8029b73",
  1590 => x"d3e8c187",
  1591 => x"d1ebc049",
  1592 => x"fadfff87",
  1593 => x"1e731e87",
  1594 => x"4bffc31e",
  1595 => x"fc4ad4ff",
  1596 => x"98c148bf",
  1597 => x"026e7e70",
  1598 => x"ff87fbc0",
  1599 => x"c1c148d0",
  1600 => x"7ad2c278",
  1601 => x"d1c37a73",
  1602 => x"ff4849c7",
  1603 => x"73506a80",
  1604 => x"73516a7a",
  1605 => x"6a80c17a",
  1606 => x"6a7a7350",
  1607 => x"6a7a7350",
  1608 => x"6a7a7349",
  1609 => x"6a7a7350",
  1610 => x"d0d1c350",
  1611 => x"d0ff5997",
  1612 => x"78c0c148",
  1613 => x"d1c387d7",
  1614 => x"ff4849c7",
  1615 => x"5150c080",
  1616 => x"50c080c1",
  1617 => x"50c150d9",
  1618 => x"c350e2c0",
  1619 => x"cdd1c350",
  1620 => x"f850c048",
  1621 => x"deff2680",
  1622 => x"c71e87c5",
  1623 => x"49c187f7",
  1624 => x"fe87c4fd",
  1625 => x"7087c6e7",
  1626 => x"87cd0298",
  1627 => x"87c3f0fe",
  1628 => x"c4029870",
  1629 => x"c24ac187",
  1630 => x"724ac087",
  1631 => x"87ce059a",
  1632 => x"e6c11ec0",
  1633 => x"f5c049ef",
  1634 => x"86c487f7",
  1635 => x"e6c187fe",
  1636 => x"1ec087ed",
  1637 => x"49fae6c1",
  1638 => x"87e5f5c0",
  1639 => x"e7c11ec0",
  1640 => x"497087c6",
  1641 => x"87d9f5c0",
  1642 => x"f887e9c3",
  1643 => x"534f268e",
  1644 => x"61662044",
  1645 => x"64656c69",
  1646 => x"6f42002e",
  1647 => x"6e69746f",
  1648 => x"2e2e2e67",
  1649 => x"c01e1e00",
  1650 => x"c187c3ec",
  1651 => x"6e87dcda",
  1652 => x"ffffc149",
  1653 => x"c1486e99",
  1654 => x"717e7080",
  1655 => x"87e70599",
  1656 => x"7087c2fc",
  1657 => x"87f5ce49",
  1658 => x"2687dcff",
  1659 => x"c31e4f26",
  1660 => x"c048fcdd",
  1661 => x"f8ddc378",
  1662 => x"fd78c048",
  1663 => x"c4ff87dc",
  1664 => x"2648c087",
  1665 => x"4520804f",
  1666 => x"00746978",
  1667 => x"61422080",
  1668 => x"21006b63",
  1669 => x"91000013",
  1670 => x"00000037",
  1671 => x"13210000",
  1672 => x"37af0000",
  1673 => x"00000000",
  1674 => x"00132100",
  1675 => x"0037cd00",
  1676 => x"00000000",
  1677 => x"00001321",
  1678 => x"000037eb",
  1679 => x"21000000",
  1680 => x"09000013",
  1681 => x"00000038",
  1682 => x"13210000",
  1683 => x"38270000",
  1684 => x"00000000",
  1685 => x"00132100",
  1686 => x"00384500",
  1687 => x"00000000",
  1688 => x"00001321",
  1689 => x"00000000",
  1690 => x"bc000000",
  1691 => x"00000013",
  1692 => x"00000000",
  1693 => x"6f4c0000",
  1694 => x"2a206461",
  1695 => x"fe1e002e",
  1696 => x"78c048f0",
  1697 => x"097909cd",
  1698 => x"1e1e4f26",
  1699 => x"7ebff0fe",
  1700 => x"4f262648",
  1701 => x"48f0fe1e",
  1702 => x"4f2678c1",
  1703 => x"48f0fe1e",
  1704 => x"4f2678c0",
  1705 => x"c04a711e",
  1706 => x"4f265252",
  1707 => x"5c5b5e0e",
  1708 => x"86f40e5d",
  1709 => x"6d974d71",
  1710 => x"4ca5c17e",
  1711 => x"c8486c97",
  1712 => x"486e58a6",
  1713 => x"05a866c4",
  1714 => x"48ff87c5",
  1715 => x"ff87e6c0",
  1716 => x"a5c287ca",
  1717 => x"4b6c9749",
  1718 => x"974ba371",
  1719 => x"6c974b6b",
  1720 => x"c1486e7e",
  1721 => x"58a6c880",
  1722 => x"a6cc98c7",
  1723 => x"7c977058",
  1724 => x"7387e1fe",
  1725 => x"268ef448",
  1726 => x"264c264d",
  1727 => x"0e4f264b",
  1728 => x"0e5c5b5e",
  1729 => x"4c7186f4",
  1730 => x"c34a66d8",
  1731 => x"a4c29aff",
  1732 => x"496c974b",
  1733 => x"7249a173",
  1734 => x"7e6c9751",
  1735 => x"80c1486e",
  1736 => x"c758a6c8",
  1737 => x"58a6cc98",
  1738 => x"8ef45470",
  1739 => x"1e87caff",
  1740 => x"87e8fd1e",
  1741 => x"494abfe0",
  1742 => x"99c0e0c0",
  1743 => x"7287cb02",
  1744 => x"e3e1c31e",
  1745 => x"87f7fe49",
  1746 => x"fdfc86c4",
  1747 => x"fd7e7087",
  1748 => x"262687c2",
  1749 => x"e1c31e4f",
  1750 => x"c7fd49e3",
  1751 => x"efecc187",
  1752 => x"87dafc49",
  1753 => x"2687d9c5",
  1754 => x"5b5e0e4f",
  1755 => x"c30e5d5c",
  1756 => x"4abfc6e2",
  1757 => x"bffdeec1",
  1758 => x"bc724c49",
  1759 => x"dbfc4d71",
  1760 => x"744bc087",
  1761 => x"0299d049",
  1762 => x"497587d5",
  1763 => x"1e7199d0",
  1764 => x"f5c11ec0",
  1765 => x"82734acf",
  1766 => x"e4c04912",
  1767 => x"c186c887",
  1768 => x"c8832d2c",
  1769 => x"daff04ab",
  1770 => x"87e8fb87",
  1771 => x"48fdeec1",
  1772 => x"bfc6e2c3",
  1773 => x"264d2678",
  1774 => x"264b264c",
  1775 => x"0000004f",
  1776 => x"d0ff1e00",
  1777 => x"78e1c848",
  1778 => x"c548d4ff",
  1779 => x"0266c478",
  1780 => x"e0c387c3",
  1781 => x"0266c878",
  1782 => x"d4ff87c6",
  1783 => x"78f0c348",
  1784 => x"7148d4ff",
  1785 => x"48d0ff78",
  1786 => x"c078e1c8",
  1787 => x"4f2678e0",
  1788 => x"5c5b5e0e",
  1789 => x"c34c710e",
  1790 => x"fa49e3e1",
  1791 => x"4a7087ee",
  1792 => x"04aab7c0",
  1793 => x"c387e3c2",
  1794 => x"c905aae0",
  1795 => x"f3f2c187",
  1796 => x"c278c148",
  1797 => x"f0c387d4",
  1798 => x"87c905aa",
  1799 => x"48eff2c1",
  1800 => x"f5c178c1",
  1801 => x"f3f2c187",
  1802 => x"87c702bf",
  1803 => x"c0c24b72",
  1804 => x"7287c2b3",
  1805 => x"059c744b",
  1806 => x"f2c187d1",
  1807 => x"c11ebfef",
  1808 => x"1ebff3f2",
  1809 => x"f8fd4972",
  1810 => x"c186c887",
  1811 => x"02bfeff2",
  1812 => x"7387e0c0",
  1813 => x"29b7c449",
  1814 => x"cff4c191",
  1815 => x"cf4a7381",
  1816 => x"c192c29a",
  1817 => x"70307248",
  1818 => x"72baff4a",
  1819 => x"70986948",
  1820 => x"7387db79",
  1821 => x"29b7c449",
  1822 => x"cff4c191",
  1823 => x"cf4a7381",
  1824 => x"c392c29a",
  1825 => x"70307248",
  1826 => x"b069484a",
  1827 => x"f2c17970",
  1828 => x"78c048f3",
  1829 => x"48eff2c1",
  1830 => x"e1c378c0",
  1831 => x"cbf849e3",
  1832 => x"c04a7087",
  1833 => x"fd03aab7",
  1834 => x"48c087dd",
  1835 => x"0087c8fc",
  1836 => x"00000000",
  1837 => x"1e000000",
  1838 => x"fc494a71",
  1839 => x"4f2687f2",
  1840 => x"724ac01e",
  1841 => x"c191c449",
  1842 => x"c081cff4",
  1843 => x"d082c179",
  1844 => x"ee04aab7",
  1845 => x"0e4f2687",
  1846 => x"5d5c5b5e",
  1847 => x"f64d710e",
  1848 => x"4a7587fa",
  1849 => x"922ab7c4",
  1850 => x"82cff4c1",
  1851 => x"9ccf4c75",
  1852 => x"496a94c2",
  1853 => x"c32b744b",
  1854 => x"7448c29b",
  1855 => x"ff4c7030",
  1856 => x"714874bc",
  1857 => x"f67a7098",
  1858 => x"487387ca",
  1859 => x"0087e6fa",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"00000000",
  1868 => x"00000000",
  1869 => x"00000000",
  1870 => x"00000000",
  1871 => x"00000000",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00000000",
  1875 => x"16000000",
  1876 => x"2e25261e",
  1877 => x"1e3e3d36",
  1878 => x"c848d0ff",
  1879 => x"487178e1",
  1880 => x"7808d4ff",
  1881 => x"ff1e4f26",
  1882 => x"e1c848d0",
  1883 => x"ff487178",
  1884 => x"c47808d4",
  1885 => x"d4ff4866",
  1886 => x"4f267808",
  1887 => x"c44a711e",
  1888 => x"e0c11e66",
  1889 => x"ddff49a2",
  1890 => x"4966c887",
  1891 => x"ff29b7c8",
  1892 => x"787148d4",
  1893 => x"c048d0ff",
  1894 => x"262678e0",
  1895 => x"1e731e4f",
  1896 => x"e2c04b71",
  1897 => x"87effe49",
  1898 => x"48134ac7",
  1899 => x"7808d4ff",
  1900 => x"8ac14972",
  1901 => x"f1059971",
  1902 => x"48d0ff87",
  1903 => x"c478e0c0",
  1904 => x"264d2687",
  1905 => x"264b264c",
  1906 => x"d4ff1e4f",
  1907 => x"7affc34a",
  1908 => x"c848d0ff",
  1909 => x"7ade78e1",
  1910 => x"bfede1c3",
  1911 => x"c848497a",
  1912 => x"717a7028",
  1913 => x"7028d048",
  1914 => x"d848717a",
  1915 => x"c37a7028",
  1916 => x"7abff1e1",
  1917 => x"28c84849",
  1918 => x"48717a70",
  1919 => x"7a7028d0",
  1920 => x"28d84871",
  1921 => x"d0ff7a70",
  1922 => x"78e0c048",
  1923 => x"731e4f26",
  1924 => x"c34a711e",
  1925 => x"4bbfede1",
  1926 => x"e0c02b72",
  1927 => x"87ce04aa",
  1928 => x"e0c04972",
  1929 => x"f1e1c389",
  1930 => x"2b714bbf",
  1931 => x"e0c087cf",
  1932 => x"c3897249",
  1933 => x"48bff1e1",
  1934 => x"49703071",
  1935 => x"9b66c8b3",
  1936 => x"87c44873",
  1937 => x"4c264d26",
  1938 => x"4f264b26",
  1939 => x"5c5b5e0e",
  1940 => x"86ec0e5d",
  1941 => x"e1c34b71",
  1942 => x"4c7ebfed",
  1943 => x"e0c02c73",
  1944 => x"e0c004ab",
  1945 => x"48a6c487",
  1946 => x"497378c0",
  1947 => x"7189e0c0",
  1948 => x"66e4c04a",
  1949 => x"cc307248",
  1950 => x"e1c358a6",
  1951 => x"4c4dbff1",
  1952 => x"e4c02c71",
  1953 => x"c0497387",
  1954 => x"714866e4",
  1955 => x"58a6c830",
  1956 => x"7349e0c0",
  1957 => x"66e4c089",
  1958 => x"cc287148",
  1959 => x"e1c358a6",
  1960 => x"484dbff1",
  1961 => x"49703071",
  1962 => x"66e4c0b4",
  1963 => x"c084c19c",
  1964 => x"04ac66e8",
  1965 => x"4cc087c2",
  1966 => x"04abe0c0",
  1967 => x"a6cc87d3",
  1968 => x"7378c048",
  1969 => x"89e0c049",
  1970 => x"30714874",
  1971 => x"d558a6d4",
  1972 => x"74497387",
  1973 => x"d0307148",
  1974 => x"e0c058a6",
  1975 => x"74897349",
  1976 => x"d4287148",
  1977 => x"66c458a6",
  1978 => x"6ebaff4a",
  1979 => x"4966c89a",
  1980 => x"9975b9ff",
  1981 => x"66cc4872",
  1982 => x"f1e1c3b0",
  1983 => x"d0487158",
  1984 => x"e1c3b066",
  1985 => x"c0fb58f5",
  1986 => x"fc8eec87",
  1987 => x"ff1e87f6",
  1988 => x"c9c848d0",
  1989 => x"ff487178",
  1990 => x"267808d4",
  1991 => x"4a711e4f",
  1992 => x"ff87eb49",
  1993 => x"78c848d0",
  1994 => x"731e4f26",
  1995 => x"c34b711e",
  1996 => x"02bfc1e2",
  1997 => x"ebc287c3",
  1998 => x"48d0ff87",
  1999 => x"7378c9c8",
  2000 => x"b1e0c049",
  2001 => x"7148d4ff",
  2002 => x"f5e1c378",
  2003 => x"c878c048",
  2004 => x"87c50266",
  2005 => x"c249ffc3",
  2006 => x"c349c087",
  2007 => x"cc59fde1",
  2008 => x"87c60266",
  2009 => x"4ad5d5c5",
  2010 => x"ffcf87c4",
  2011 => x"e2c34aff",
  2012 => x"e2c35ac1",
  2013 => x"78c148c1",
  2014 => x"4d2687c4",
  2015 => x"4b264c26",
  2016 => x"5e0e4f26",
  2017 => x"0e5d5c5b",
  2018 => x"e1c34a71",
  2019 => x"724cbffd",
  2020 => x"87cb029a",
  2021 => x"c191c849",
  2022 => x"714be0fc",
  2023 => x"c287c483",
  2024 => x"c04be0c0",
  2025 => x"7449134d",
  2026 => x"f9e1c399",
  2027 => x"d4ffb9bf",
  2028 => x"c1787148",
  2029 => x"c8852cb7",
  2030 => x"e804adb7",
  2031 => x"f5e1c387",
  2032 => x"80c848bf",
  2033 => x"58f9e1c3",
  2034 => x"1e87effe",
  2035 => x"4b711e73",
  2036 => x"029a4a13",
  2037 => x"497287cb",
  2038 => x"1387e7fe",
  2039 => x"f5059a4a",
  2040 => x"87dafe87",
  2041 => x"f5e1c31e",
  2042 => x"e1c349bf",
  2043 => x"a1c148f5",
  2044 => x"b7c0c478",
  2045 => x"87db03a9",
  2046 => x"c348d4ff",
  2047 => x"78bff9e1",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
