library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4eac387",
    12 => x"86c0c64e",
    13 => x"49c4eac3",
    14 => x"48e0d0c3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e3e6",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"731e4f26",
    53 => x"029a721e",
    54 => x"c087e7c0",
    55 => x"724bc148",
    56 => x"87d106a9",
    57 => x"c9068272",
    58 => x"72837387",
    59 => x"87f401a9",
    60 => x"b2c187c3",
    61 => x"03a9723a",
    62 => x"07807389",
    63 => x"052b2ac1",
    64 => x"4b2687f3",
    65 => x"751e4f26",
    66 => x"714dc41e",
    67 => x"ff04a1b7",
    68 => x"c381c1b9",
    69 => x"b77207bd",
    70 => x"baff04a2",
    71 => x"bdc182c1",
    72 => x"87eefe07",
    73 => x"ff042dc1",
    74 => x"0780c1b8",
    75 => x"b9ff042d",
    76 => x"260781c1",
    77 => x"1e4f264d",
    78 => x"d4ff4811",
    79 => x"66c47808",
    80 => x"c888c148",
    81 => x"987058a6",
    82 => x"2687ed05",
    83 => x"d4ff1e4f",
    84 => x"78ffc348",
    85 => x"66c45168",
    86 => x"c888c148",
    87 => x"987058a6",
    88 => x"2687eb05",
    89 => x"1e731e4f",
    90 => x"c34bd4ff",
    91 => x"4a6b7bff",
    92 => x"6b7bffc3",
    93 => x"7232c849",
    94 => x"7bffc3b1",
    95 => x"31c84a6b",
    96 => x"ffc3b271",
    97 => x"c8496b7b",
    98 => x"71b17232",
    99 => x"2687c448",
   100 => x"264c264d",
   101 => x"0e4f264b",
   102 => x"5d5c5b5e",
   103 => x"ff4a710e",
   104 => x"49724cd4",
   105 => x"7199ffc3",
   106 => x"e0d0c37c",
   107 => x"87c805bf",
   108 => x"c94866d0",
   109 => x"58a6d430",
   110 => x"d84966d0",
   111 => x"99ffc329",
   112 => x"66d07c71",
   113 => x"c329d049",
   114 => x"7c7199ff",
   115 => x"c84966d0",
   116 => x"99ffc329",
   117 => x"66d07c71",
   118 => x"99ffc349",
   119 => x"49727c71",
   120 => x"ffc329d0",
   121 => x"6c7c7199",
   122 => x"fff0c94b",
   123 => x"abffc34d",
   124 => x"c387d005",
   125 => x"4b6c7cff",
   126 => x"c6028dc1",
   127 => x"abffc387",
   128 => x"7387f002",
   129 => x"87c7fe48",
   130 => x"ff49c01e",
   131 => x"ffc348d4",
   132 => x"c381c178",
   133 => x"04a9b7c8",
   134 => x"4f2687f1",
   135 => x"e71e731e",
   136 => x"dff8c487",
   137 => x"c01ec04b",
   138 => x"f7c1f0ff",
   139 => x"87e7fd49",
   140 => x"a8c186c4",
   141 => x"87eac005",
   142 => x"c348d4ff",
   143 => x"c0c178ff",
   144 => x"c0c0c0c0",
   145 => x"f0e1c01e",
   146 => x"fd49e9c1",
   147 => x"86c487c9",
   148 => x"ca059870",
   149 => x"48d4ff87",
   150 => x"c178ffc3",
   151 => x"fe87cb48",
   152 => x"8bc187e6",
   153 => x"87fdfe05",
   154 => x"e6fc48c0",
   155 => x"1e731e87",
   156 => x"c348d4ff",
   157 => x"4bd378ff",
   158 => x"ffc01ec0",
   159 => x"49c1c1f0",
   160 => x"c487d4fc",
   161 => x"05987086",
   162 => x"d4ff87ca",
   163 => x"78ffc348",
   164 => x"87cb48c1",
   165 => x"c187f1fd",
   166 => x"dbff058b",
   167 => x"fb48c087",
   168 => x"5e0e87f1",
   169 => x"ff0e5c5b",
   170 => x"dbfd4cd4",
   171 => x"1eeac687",
   172 => x"c1f0e1c0",
   173 => x"defb49c8",
   174 => x"c186c487",
   175 => x"87c802a8",
   176 => x"c087eafe",
   177 => x"87e2c148",
   178 => x"7087dafa",
   179 => x"ffffcf49",
   180 => x"a9eac699",
   181 => x"fe87c802",
   182 => x"48c087d3",
   183 => x"c387cbc1",
   184 => x"f1c07cff",
   185 => x"87f4fc4b",
   186 => x"c0029870",
   187 => x"1ec087eb",
   188 => x"c1f0ffc0",
   189 => x"defa49fa",
   190 => x"7086c487",
   191 => x"87d90598",
   192 => x"6c7cffc3",
   193 => x"7cffc349",
   194 => x"c17c7c7c",
   195 => x"c40299c0",
   196 => x"d548c187",
   197 => x"d148c087",
   198 => x"05abc287",
   199 => x"48c087c4",
   200 => x"8bc187c8",
   201 => x"87fdfe05",
   202 => x"e4f948c0",
   203 => x"1e731e87",
   204 => x"48e0d0c3",
   205 => x"4bc778c1",
   206 => x"c248d0ff",
   207 => x"87c8fb78",
   208 => x"c348d0ff",
   209 => x"c01ec078",
   210 => x"c0c1d0e5",
   211 => x"87c7f949",
   212 => x"a8c186c4",
   213 => x"4b87c105",
   214 => x"c505abc2",
   215 => x"c048c087",
   216 => x"8bc187f9",
   217 => x"87d0ff05",
   218 => x"c387f7fc",
   219 => x"7058e4d0",
   220 => x"87cd0598",
   221 => x"ffc01ec1",
   222 => x"49d0c1f0",
   223 => x"c487d8f8",
   224 => x"48d4ff86",
   225 => x"c478ffc3",
   226 => x"d0c387e0",
   227 => x"d0ff58e8",
   228 => x"ff78c248",
   229 => x"ffc348d4",
   230 => x"f748c178",
   231 => x"5e0e87f5",
   232 => x"0e5d5c5b",
   233 => x"ffc34a71",
   234 => x"4cd4ff4d",
   235 => x"d0ff7c75",
   236 => x"78c3c448",
   237 => x"1e727c75",
   238 => x"c1f0ffc0",
   239 => x"d6f749d8",
   240 => x"7086c487",
   241 => x"87c50298",
   242 => x"f0c048c0",
   243 => x"c37c7587",
   244 => x"c0c87cfe",
   245 => x"4966d41e",
   246 => x"c487dcf5",
   247 => x"757c7586",
   248 => x"d87c757c",
   249 => x"754be0da",
   250 => x"99496c7c",
   251 => x"c187c505",
   252 => x"87f3058b",
   253 => x"d0ff7c75",
   254 => x"c178c248",
   255 => x"87cff648",
   256 => x"4ad4ff1e",
   257 => x"c448d0ff",
   258 => x"ffc378d1",
   259 => x"0589c17a",
   260 => x"4f2687f8",
   261 => x"711e731e",
   262 => x"cdeec54b",
   263 => x"d4ff4adf",
   264 => x"78ffc348",
   265 => x"fec34868",
   266 => x"87c502a8",
   267 => x"ed058ac1",
   268 => x"059a7287",
   269 => x"48c087c5",
   270 => x"7387eac0",
   271 => x"87cc029b",
   272 => x"731e66c8",
   273 => x"87c5f449",
   274 => x"87c686c4",
   275 => x"fe4966c8",
   276 => x"d4ff87ee",
   277 => x"78ffc348",
   278 => x"059b7378",
   279 => x"d0ff87c5",
   280 => x"c178d048",
   281 => x"87ebf448",
   282 => x"711e731e",
   283 => x"ff4bc04a",
   284 => x"ffc348d4",
   285 => x"48d0ff78",
   286 => x"ff78c3c4",
   287 => x"ffc348d4",
   288 => x"c01e7278",
   289 => x"d1c1f0ff",
   290 => x"87cbf449",
   291 => x"987086c4",
   292 => x"c887cd05",
   293 => x"66cc1ec0",
   294 => x"87f8fd49",
   295 => x"4b7086c4",
   296 => x"c248d0ff",
   297 => x"f3487378",
   298 => x"5e0e87e9",
   299 => x"0e5d5c5b",
   300 => x"ffc01ec0",
   301 => x"49c9c1f0",
   302 => x"d287dcf3",
   303 => x"e8d0c31e",
   304 => x"87d0fd49",
   305 => x"4cc086c8",
   306 => x"b7d284c1",
   307 => x"87f804ac",
   308 => x"97e8d0c3",
   309 => x"c0c349bf",
   310 => x"a9c0c199",
   311 => x"87e7c005",
   312 => x"97efd0c3",
   313 => x"31d049bf",
   314 => x"97f0d0c3",
   315 => x"32c84abf",
   316 => x"d0c3b172",
   317 => x"4abf97f1",
   318 => x"cf4c71b1",
   319 => x"9cffffff",
   320 => x"34ca84c1",
   321 => x"c387e7c1",
   322 => x"bf97f1d0",
   323 => x"c631c149",
   324 => x"f2d0c399",
   325 => x"c74abf97",
   326 => x"b1722ab7",
   327 => x"97edd0c3",
   328 => x"cf4d4abf",
   329 => x"eed0c39d",
   330 => x"c34abf97",
   331 => x"c332ca9a",
   332 => x"bf97efd0",
   333 => x"7333c24b",
   334 => x"f0d0c3b2",
   335 => x"c34bbf97",
   336 => x"b7c69bc0",
   337 => x"c2b2732b",
   338 => x"7148c181",
   339 => x"c1497030",
   340 => x"70307548",
   341 => x"c14c724d",
   342 => x"c8947184",
   343 => x"06adb7c0",
   344 => x"34c187cc",
   345 => x"c0c82db7",
   346 => x"ff01adb7",
   347 => x"487487f4",
   348 => x"0e87dcf0",
   349 => x"5d5c5b5e",
   350 => x"c386f80e",
   351 => x"c048ced9",
   352 => x"c6d1c378",
   353 => x"fb49c01e",
   354 => x"86c487de",
   355 => x"c5059870",
   356 => x"c948c087",
   357 => x"4dc087ce",
   358 => x"fac07ec1",
   359 => x"c349bff2",
   360 => x"714afcd1",
   361 => x"c1eb4bc8",
   362 => x"05987087",
   363 => x"7ec087c2",
   364 => x"bfeefac0",
   365 => x"d8d2c349",
   366 => x"4bc8714a",
   367 => x"7087ebea",
   368 => x"87c20598",
   369 => x"026e7ec0",
   370 => x"c387fdc0",
   371 => x"4dbfccd8",
   372 => x"9fc4d9c3",
   373 => x"c5487ebf",
   374 => x"05a8ead6",
   375 => x"d8c387c7",
   376 => x"ce4dbfcc",
   377 => x"ca486e87",
   378 => x"02a8d5e9",
   379 => x"48c087c5",
   380 => x"c387f1c7",
   381 => x"751ec6d1",
   382 => x"87ecf949",
   383 => x"987086c4",
   384 => x"c087c505",
   385 => x"87dcc748",
   386 => x"bfeefac0",
   387 => x"d8d2c349",
   388 => x"4bc8714a",
   389 => x"7087d3e9",
   390 => x"87c80598",
   391 => x"48ced9c3",
   392 => x"87da78c1",
   393 => x"bff2fac0",
   394 => x"fcd1c349",
   395 => x"4bc8714a",
   396 => x"7087f7e8",
   397 => x"c5c00298",
   398 => x"c648c087",
   399 => x"d9c387e6",
   400 => x"49bf97c4",
   401 => x"05a9d5c1",
   402 => x"c387cdc0",
   403 => x"bf97c5d9",
   404 => x"a9eac249",
   405 => x"87c5c002",
   406 => x"c7c648c0",
   407 => x"c6d1c387",
   408 => x"487ebf97",
   409 => x"02a8e9c3",
   410 => x"6e87cec0",
   411 => x"a8ebc348",
   412 => x"87c5c002",
   413 => x"ebc548c0",
   414 => x"d1d1c387",
   415 => x"9949bf97",
   416 => x"87ccc005",
   417 => x"97d2d1c3",
   418 => x"a9c249bf",
   419 => x"87c5c002",
   420 => x"cfc548c0",
   421 => x"d3d1c387",
   422 => x"c348bf97",
   423 => x"7058cad9",
   424 => x"88c1484c",
   425 => x"58ced9c3",
   426 => x"97d4d1c3",
   427 => x"817549bf",
   428 => x"97d5d1c3",
   429 => x"32c84abf",
   430 => x"c37ea172",
   431 => x"6e48dbdd",
   432 => x"d6d1c378",
   433 => x"c848bf97",
   434 => x"d9c358a6",
   435 => x"c202bfce",
   436 => x"fac087d4",
   437 => x"c349bfee",
   438 => x"714ad8d2",
   439 => x"c9e64bc8",
   440 => x"02987087",
   441 => x"c087c5c0",
   442 => x"87f8c348",
   443 => x"bfc6d9c3",
   444 => x"efddc34c",
   445 => x"ebd1c35c",
   446 => x"c849bf97",
   447 => x"ead1c331",
   448 => x"a14abf97",
   449 => x"ecd1c349",
   450 => x"d04abf97",
   451 => x"49a17232",
   452 => x"97edd1c3",
   453 => x"32d84abf",
   454 => x"c449a172",
   455 => x"ddc39166",
   456 => x"c381bfdb",
   457 => x"c359e3dd",
   458 => x"bf97f3d1",
   459 => x"c332c84a",
   460 => x"bf97f2d1",
   461 => x"c34aa24b",
   462 => x"bf97f4d1",
   463 => x"7333d04b",
   464 => x"d1c34aa2",
   465 => x"4bbf97f5",
   466 => x"33d89bcf",
   467 => x"c34aa273",
   468 => x"c35ae7dd",
   469 => x"4abfe3dd",
   470 => x"92748ac2",
   471 => x"48e7ddc3",
   472 => x"c178a172",
   473 => x"d1c387ca",
   474 => x"49bf97d8",
   475 => x"d1c331c8",
   476 => x"4abf97d7",
   477 => x"d9c349a1",
   478 => x"d9c359d6",
   479 => x"c549bfd2",
   480 => x"81ffc731",
   481 => x"ddc329c9",
   482 => x"d1c359ef",
   483 => x"4abf97dd",
   484 => x"d1c332c8",
   485 => x"4bbf97dc",
   486 => x"66c44aa2",
   487 => x"c3826e92",
   488 => x"c35aebdd",
   489 => x"c048e3dd",
   490 => x"dfddc378",
   491 => x"78a17248",
   492 => x"48efddc3",
   493 => x"bfe3ddc3",
   494 => x"f3ddc378",
   495 => x"e7ddc348",
   496 => x"d9c378bf",
   497 => x"c002bfce",
   498 => x"487487c9",
   499 => x"7e7030c4",
   500 => x"c387c9c0",
   501 => x"48bfebdd",
   502 => x"7e7030c4",
   503 => x"48d2d9c3",
   504 => x"48c1786e",
   505 => x"4d268ef8",
   506 => x"4b264c26",
   507 => x"5e0e4f26",
   508 => x"0e5d5c5b",
   509 => x"d9c34a71",
   510 => x"cb02bfce",
   511 => x"c74b7287",
   512 => x"c14c722b",
   513 => x"87c99cff",
   514 => x"2bc84b72",
   515 => x"ffc34c72",
   516 => x"dbddc39c",
   517 => x"fac083bf",
   518 => x"02abbfea",
   519 => x"fac087d9",
   520 => x"d1c35bee",
   521 => x"49731ec6",
   522 => x"c487fdf0",
   523 => x"05987086",
   524 => x"48c087c5",
   525 => x"c387e6c0",
   526 => x"02bfced9",
   527 => x"497487d2",
   528 => x"d1c391c4",
   529 => x"4d6981c6",
   530 => x"ffffffcf",
   531 => x"87cb9dff",
   532 => x"91c24974",
   533 => x"81c6d1c3",
   534 => x"754d699f",
   535 => x"87c6fe48",
   536 => x"5c5b5e0e",
   537 => x"711e0e5d",
   538 => x"c11ec04d",
   539 => x"87e2d149",
   540 => x"4c7086c4",
   541 => x"c2c1029c",
   542 => x"d6d9c387",
   543 => x"ff49754a",
   544 => x"7087ccdf",
   545 => x"f2c00298",
   546 => x"754a7487",
   547 => x"ff4bcb49",
   548 => x"7087f1df",
   549 => x"e2c00298",
   550 => x"741ec087",
   551 => x"87c7029c",
   552 => x"c048a6c4",
   553 => x"c487c578",
   554 => x"78c148a6",
   555 => x"d04966c4",
   556 => x"86c487e0",
   557 => x"059c4c70",
   558 => x"7487fefe",
   559 => x"e5fc2648",
   560 => x"5b5e0e87",
   561 => x"f80e5d5c",
   562 => x"9b4b7186",
   563 => x"c087c505",
   564 => x"87d4c248",
   565 => x"c04da3c8",
   566 => x"0266d87d",
   567 => x"66d887c7",
   568 => x"c505bf97",
   569 => x"c148c087",
   570 => x"66d887fe",
   571 => x"87f0fd49",
   572 => x"026e7e70",
   573 => x"6e87efc1",
   574 => x"6981dc49",
   575 => x"da496e7d",
   576 => x"4ca3c481",
   577 => x"c37c699f",
   578 => x"02bfced9",
   579 => x"496e87d0",
   580 => x"699f81d4",
   581 => x"ffc04a49",
   582 => x"32d09aff",
   583 => x"4ac087c2",
   584 => x"6c484972",
   585 => x"c07c7080",
   586 => x"49a3cc7b",
   587 => x"a3d0796c",
   588 => x"c479c049",
   589 => x"78c048a6",
   590 => x"c44aa3d4",
   591 => x"91c84966",
   592 => x"c049a172",
   593 => x"c4796c41",
   594 => x"80c14866",
   595 => x"d058a6c8",
   596 => x"ff04a8b7",
   597 => x"4a6d87e2",
   598 => x"2ac72ac9",
   599 => x"49a3d4c2",
   600 => x"486e7972",
   601 => x"48c087c2",
   602 => x"f9f98ef8",
   603 => x"5b5e0e87",
   604 => x"710e5d5c",
   605 => x"eafac04c",
   606 => x"7478ff48",
   607 => x"cac1029c",
   608 => x"49a4c887",
   609 => x"c2c10269",
   610 => x"4a66d087",
   611 => x"d482496c",
   612 => x"66d05aa6",
   613 => x"d9c3b94d",
   614 => x"ff4abfca",
   615 => x"719972ba",
   616 => x"e4c00299",
   617 => x"4ba4c487",
   618 => x"c1f9496b",
   619 => x"c37b7087",
   620 => x"49bfc6d9",
   621 => x"7c71816c",
   622 => x"d9c3b975",
   623 => x"ff4abfca",
   624 => x"719972ba",
   625 => x"dcff0599",
   626 => x"f87c7587",
   627 => x"731e87d8",
   628 => x"9b4b711e",
   629 => x"c887c702",
   630 => x"056949a3",
   631 => x"48c087c5",
   632 => x"c387ebc0",
   633 => x"4abfdfdd",
   634 => x"6949a3c4",
   635 => x"c389c249",
   636 => x"91bfc6d9",
   637 => x"c34aa271",
   638 => x"49bfcad9",
   639 => x"a271996b",
   640 => x"1e66c84a",
   641 => x"dfe94972",
   642 => x"7086c487",
   643 => x"d9f74849",
   644 => x"1e731e87",
   645 => x"029b4b71",
   646 => x"a3c887c7",
   647 => x"c5056949",
   648 => x"c048c087",
   649 => x"ddc387eb",
   650 => x"c44abfdf",
   651 => x"496949a3",
   652 => x"d9c389c2",
   653 => x"7191bfc6",
   654 => x"d9c34aa2",
   655 => x"6b49bfca",
   656 => x"4aa27199",
   657 => x"721e66c8",
   658 => x"87d2e549",
   659 => x"497086c4",
   660 => x"87d6f648",
   661 => x"5c5b5e0e",
   662 => x"86f80e5d",
   663 => x"a6c44b71",
   664 => x"c878ff48",
   665 => x"4d6949a3",
   666 => x"a3d44cc0",
   667 => x"c849744a",
   668 => x"49a17291",
   669 => x"66d84969",
   670 => x"70887148",
   671 => x"a966d87e",
   672 => x"6e87ca01",
   673 => x"87c506ad",
   674 => x"6e5ca6c8",
   675 => x"d084c14d",
   676 => x"ff04acb7",
   677 => x"66c487d4",
   678 => x"f58ef848",
   679 => x"5e0e87c8",
   680 => x"0e5d5c5b",
   681 => x"a6c886ec",
   682 => x"48a6c859",
   683 => x"ffffffc1",
   684 => x"c478ffff",
   685 => x"c078ff80",
   686 => x"c44cc04d",
   687 => x"83d44b66",
   688 => x"91c84974",
   689 => x"7549a173",
   690 => x"7392c84a",
   691 => x"49697ea2",
   692 => x"d489bf6e",
   693 => x"ad7459a6",
   694 => x"d087c605",
   695 => x"bf6e48a6",
   696 => x"4866d078",
   697 => x"04a8b7c0",
   698 => x"66d087cf",
   699 => x"a966c849",
   700 => x"d087c603",
   701 => x"a6cc5ca6",
   702 => x"d084c159",
   703 => x"fe04acb7",
   704 => x"85c187f9",
   705 => x"04adb7d0",
   706 => x"cc87eefe",
   707 => x"8eec4866",
   708 => x"0e87d3f3",
   709 => x"0e5c5b5e",
   710 => x"4cc04b71",
   711 => x"6949a3c8",
   712 => x"7429c449",
   713 => x"1e71914a",
   714 => x"87d44973",
   715 => x"84c186c4",
   716 => x"04acb7d0",
   717 => x"1ec087e6",
   718 => x"87c44973",
   719 => x"87e8f226",
   720 => x"5c5b5e0e",
   721 => x"86f00e5d",
   722 => x"e0c04b71",
   723 => x"2cc94c66",
   724 => x"c3029b73",
   725 => x"a3c887e1",
   726 => x"c3026949",
   727 => x"a3d087d9",
   728 => x"66e0c049",
   729 => x"ac7e6b79",
   730 => x"87cbc302",
   731 => x"bfcad9c3",
   732 => x"71b9ff49",
   733 => x"719a744a",
   734 => x"cc986e48",
   735 => x"a3c458a6",
   736 => x"48a6c44d",
   737 => x"66c8786d",
   738 => x"87c505aa",
   739 => x"d1c27b74",
   740 => x"731e7287",
   741 => x"87fcfa49",
   742 => x"7e7086c4",
   743 => x"a8b7c048",
   744 => x"d487d004",
   745 => x"496e4aa3",
   746 => x"a17291c8",
   747 => x"697b2149",
   748 => x"c087c77d",
   749 => x"49a3cc7b",
   750 => x"66c87d69",
   751 => x"fa49731e",
   752 => x"86c487d2",
   753 => x"d4c27e70",
   754 => x"a6cc49a3",
   755 => x"c8786948",
   756 => x"66cc4866",
   757 => x"87c906a8",
   758 => x"b7c0486e",
   759 => x"e0c004a8",
   760 => x"c0486e87",
   761 => x"c004a8b7",
   762 => x"a3d487ec",
   763 => x"c8496e4a",
   764 => x"49a17291",
   765 => x"694866c8",
   766 => x"cc497088",
   767 => x"d506a966",
   768 => x"fa497387",
   769 => x"497087d8",
   770 => x"c84aa3d4",
   771 => x"49a17291",
   772 => x"c44166c8",
   773 => x"8c6b7966",
   774 => x"731e4974",
   775 => x"87cdf549",
   776 => x"e0c086c4",
   777 => x"ffc74966",
   778 => x"87cb0299",
   779 => x"1ec6d1c3",
   780 => x"d9f64973",
   781 => x"f086c487",
   782 => x"87eaee8e",
   783 => x"711e731e",
   784 => x"c0029b4b",
   785 => x"ddc387e4",
   786 => x"4a735bf3",
   787 => x"d9c38ac2",
   788 => x"9249bfc6",
   789 => x"bfdfddc3",
   790 => x"c3807248",
   791 => x"7158f7dd",
   792 => x"c330c448",
   793 => x"c058d6d9",
   794 => x"ddc387ed",
   795 => x"ddc348ef",
   796 => x"c378bfe3",
   797 => x"c348f3dd",
   798 => x"78bfe7dd",
   799 => x"bfced9c3",
   800 => x"c387c902",
   801 => x"49bfc6d9",
   802 => x"87c731c4",
   803 => x"bfebddc3",
   804 => x"c331c449",
   805 => x"ed59d6d9",
   806 => x"5e0e87d0",
   807 => x"710e5c5b",
   808 => x"724bc04a",
   809 => x"e1c0029a",
   810 => x"49a2da87",
   811 => x"c34b699f",
   812 => x"02bfced9",
   813 => x"a2d487cf",
   814 => x"49699f49",
   815 => x"ffffc04c",
   816 => x"c234d09c",
   817 => x"744cc087",
   818 => x"4973b349",
   819 => x"ec87edfd",
   820 => x"5e0e87d6",
   821 => x"0e5d5c5b",
   822 => x"4a7186f4",
   823 => x"9a727ec0",
   824 => x"c387d802",
   825 => x"c048c2d1",
   826 => x"fad0c378",
   827 => x"f3ddc348",
   828 => x"d0c378bf",
   829 => x"ddc348fe",
   830 => x"c378bfef",
   831 => x"c048e3d9",
   832 => x"d2d9c350",
   833 => x"d1c349bf",
   834 => x"714abfc2",
   835 => x"c0c403aa",
   836 => x"cf497287",
   837 => x"e1c00599",
   838 => x"c6d1c387",
   839 => x"fad0c31e",
   840 => x"d0c349bf",
   841 => x"a1c148fa",
   842 => x"dcff7178",
   843 => x"86c487fa",
   844 => x"48e6fac0",
   845 => x"78c6d1c3",
   846 => x"fac087cc",
   847 => x"c048bfe6",
   848 => x"fac080e0",
   849 => x"d1c358ea",
   850 => x"c148bfc2",
   851 => x"c6d1c380",
   852 => x"0ea62758",
   853 => x"97bf0000",
   854 => x"029d4dbf",
   855 => x"c387e2c2",
   856 => x"c202ade5",
   857 => x"fac087db",
   858 => x"cb4bbfe6",
   859 => x"4c1149a3",
   860 => x"c105accf",
   861 => x"497587d2",
   862 => x"89c199df",
   863 => x"d9c391cd",
   864 => x"a3c181d6",
   865 => x"c351124a",
   866 => x"51124aa3",
   867 => x"124aa3c5",
   868 => x"4aa3c751",
   869 => x"a3c95112",
   870 => x"ce51124a",
   871 => x"51124aa3",
   872 => x"124aa3d0",
   873 => x"4aa3d251",
   874 => x"a3d45112",
   875 => x"d651124a",
   876 => x"51124aa3",
   877 => x"124aa3d8",
   878 => x"4aa3dc51",
   879 => x"a3de5112",
   880 => x"c151124a",
   881 => x"87f9c07e",
   882 => x"99c84974",
   883 => x"87eac005",
   884 => x"99d04974",
   885 => x"dc87d005",
   886 => x"cac00266",
   887 => x"dc497387",
   888 => x"98700f66",
   889 => x"6e87d302",
   890 => x"87c6c005",
   891 => x"48d6d9c3",
   892 => x"fac050c0",
   893 => x"c248bfe6",
   894 => x"d9c387e7",
   895 => x"50c048e3",
   896 => x"d2d9c37e",
   897 => x"d1c349bf",
   898 => x"714abfc2",
   899 => x"c0fc04aa",
   900 => x"f3ddc387",
   901 => x"c8c005bf",
   902 => x"ced9c387",
   903 => x"fec102bf",
   904 => x"eafac087",
   905 => x"c378ff48",
   906 => x"49bffed0",
   907 => x"7087ffe6",
   908 => x"c2d1c349",
   909 => x"48a6c459",
   910 => x"bffed0c3",
   911 => x"ced9c378",
   912 => x"d8c002bf",
   913 => x"4966c487",
   914 => x"ffffffcf",
   915 => x"02a999f8",
   916 => x"c087c5c0",
   917 => x"87e1c04d",
   918 => x"dcc04dc1",
   919 => x"4966c487",
   920 => x"99f8ffcf",
   921 => x"c8c002a9",
   922 => x"48a6c887",
   923 => x"c5c078c0",
   924 => x"48a6c887",
   925 => x"66c878c1",
   926 => x"059d754d",
   927 => x"c487e0c0",
   928 => x"89c24966",
   929 => x"bfc6d9c3",
   930 => x"ddc3914a",
   931 => x"c34abfdf",
   932 => x"7248fad0",
   933 => x"d1c378a1",
   934 => x"78c048c2",
   935 => x"c087e2f9",
   936 => x"e58ef448",
   937 => x"000087c0",
   938 => x"ffff0000",
   939 => x"0eb6ffff",
   940 => x"0ebf0000",
   941 => x"41460000",
   942 => x"20323354",
   943 => x"46002020",
   944 => x"36315441",
   945 => x"00202020",
   946 => x"48d4ff1e",
   947 => x"6878ffc3",
   948 => x"1e4f2648",
   949 => x"c348d4ff",
   950 => x"d0ff78ff",
   951 => x"78e1c848",
   952 => x"d448d4ff",
   953 => x"f7ddc378",
   954 => x"bfd4ff48",
   955 => x"1e4f2650",
   956 => x"c048d0ff",
   957 => x"4f2678e0",
   958 => x"87ccff1e",
   959 => x"02994970",
   960 => x"fbc087c6",
   961 => x"87f105a9",
   962 => x"4f264871",
   963 => x"5c5b5e0e",
   964 => x"c04b710e",
   965 => x"87f0fe4c",
   966 => x"02994970",
   967 => x"c087f9c0",
   968 => x"c002a9ec",
   969 => x"fbc087f2",
   970 => x"ebc002a9",
   971 => x"b766cc87",
   972 => x"87c703ac",
   973 => x"c20266d0",
   974 => x"71537187",
   975 => x"87c20299",
   976 => x"c3fe84c1",
   977 => x"99497087",
   978 => x"c087cd02",
   979 => x"c702a9ec",
   980 => x"a9fbc087",
   981 => x"87d5ff05",
   982 => x"c30266d0",
   983 => x"7b97c087",
   984 => x"05a9ecc0",
   985 => x"4a7487c4",
   986 => x"4a7487c5",
   987 => x"728a0ac0",
   988 => x"2687c248",
   989 => x"264c264d",
   990 => x"1e4f264b",
   991 => x"7087c9fd",
   992 => x"b7f0c049",
   993 => x"87ca04a9",
   994 => x"a9b7f9c0",
   995 => x"c087c301",
   996 => x"c1c189f0",
   997 => x"ca04a9b7",
   998 => x"b7dac187",
   999 => x"87c301a9",
  1000 => x"c189f7c0",
  1001 => x"04a9b7e1",
  1002 => x"fac187ca",
  1003 => x"c301a9b7",
  1004 => x"89fdc087",
  1005 => x"4f264871",
  1006 => x"5c5b5e0e",
  1007 => x"ff4a710e",
  1008 => x"49724cd4",
  1009 => x"7087eac0",
  1010 => x"c2029b4b",
  1011 => x"ff8bc187",
  1012 => x"c5c848d0",
  1013 => x"7cd5c178",
  1014 => x"31c64973",
  1015 => x"97d5ccc3",
  1016 => x"71484abf",
  1017 => x"ff7c70b0",
  1018 => x"78c448d0",
  1019 => x"c4fe4873",
  1020 => x"5b5e0e87",
  1021 => x"f80e5d5c",
  1022 => x"c04c7186",
  1023 => x"87d3fb7e",
  1024 => x"c2c14bc0",
  1025 => x"49bf97de",
  1026 => x"cf04a9c0",
  1027 => x"87e8fb87",
  1028 => x"c2c183c1",
  1029 => x"49bf97de",
  1030 => x"87f106ab",
  1031 => x"97dec2c1",
  1032 => x"87cf02bf",
  1033 => x"7087e1fa",
  1034 => x"c6029949",
  1035 => x"a9ecc087",
  1036 => x"c087f105",
  1037 => x"87d0fa4b",
  1038 => x"cbfa4d70",
  1039 => x"58a6c887",
  1040 => x"7087c5fa",
  1041 => x"c883c14a",
  1042 => x"699749a4",
  1043 => x"c702ad49",
  1044 => x"adffc087",
  1045 => x"87e7c005",
  1046 => x"9749a4c9",
  1047 => x"66c44969",
  1048 => x"87c702a9",
  1049 => x"a8ffc048",
  1050 => x"ca87d405",
  1051 => x"699749a4",
  1052 => x"c602aa49",
  1053 => x"aaffc087",
  1054 => x"c187c405",
  1055 => x"c087d07e",
  1056 => x"c602adec",
  1057 => x"adfbc087",
  1058 => x"c087c405",
  1059 => x"6e7ec14b",
  1060 => x"87e1fe02",
  1061 => x"7387d8f9",
  1062 => x"fb8ef848",
  1063 => x"0e0087d5",
  1064 => x"5d5c5b5e",
  1065 => x"4b711e0e",
  1066 => x"ab4d4cc0",
  1067 => x"87e8c004",
  1068 => x"1ef1ffc0",
  1069 => x"c4029d75",
  1070 => x"c24ac087",
  1071 => x"724ac187",
  1072 => x"87cef049",
  1073 => x"7e7086c4",
  1074 => x"056e84c1",
  1075 => x"4c7387c2",
  1076 => x"ac7385c1",
  1077 => x"87d8ff06",
  1078 => x"2626486e",
  1079 => x"264c264d",
  1080 => x"0e4f264b",
  1081 => x"5d5c5b5e",
  1082 => x"4c711e0e",
  1083 => x"c391de49",
  1084 => x"714dd1de",
  1085 => x"026d9785",
  1086 => x"c387ddc1",
  1087 => x"4abffcdd",
  1088 => x"49728274",
  1089 => x"7087d8fe",
  1090 => x"c0026e7e",
  1091 => x"dec387f3",
  1092 => x"4a6e4bc4",
  1093 => x"fefe49cb",
  1094 => x"4b7487ce",
  1095 => x"e8c193cb",
  1096 => x"83c483d3",
  1097 => x"7bdcc5c1",
  1098 => x"c8c14974",
  1099 => x"7b7587f2",
  1100 => x"97d0dec3",
  1101 => x"c31e49bf",
  1102 => x"c249c4de",
  1103 => x"c487dfc6",
  1104 => x"c1497486",
  1105 => x"c087d9c8",
  1106 => x"f8c9c149",
  1107 => x"f8ddc387",
  1108 => x"c178c048",
  1109 => x"87cfdd49",
  1110 => x"87fffd26",
  1111 => x"64616f4c",
  1112 => x"2e676e69",
  1113 => x"0e002e2e",
  1114 => x"0e5c5b5e",
  1115 => x"c34a4b71",
  1116 => x"82bffcdd",
  1117 => x"e6fc4972",
  1118 => x"9c4c7087",
  1119 => x"4987c402",
  1120 => x"c387d7ec",
  1121 => x"c048fcdd",
  1122 => x"dc49c178",
  1123 => x"ccfd87d9",
  1124 => x"5b5e0e87",
  1125 => x"f40e5d5c",
  1126 => x"c6d1c386",
  1127 => x"c44cc04d",
  1128 => x"78c048a6",
  1129 => x"bffcddc3",
  1130 => x"06a9c049",
  1131 => x"c387c1c1",
  1132 => x"9848c6d1",
  1133 => x"87f8c002",
  1134 => x"1ef1ffc0",
  1135 => x"c70266c8",
  1136 => x"48a6c487",
  1137 => x"87c578c0",
  1138 => x"c148a6c4",
  1139 => x"4966c478",
  1140 => x"c487ffeb",
  1141 => x"c14d7086",
  1142 => x"4866c484",
  1143 => x"a6c880c1",
  1144 => x"fcddc358",
  1145 => x"03ac49bf",
  1146 => x"9d7587c6",
  1147 => x"87c8ff05",
  1148 => x"9d754cc0",
  1149 => x"87e0c302",
  1150 => x"1ef1ffc0",
  1151 => x"c70266c8",
  1152 => x"48a6cc87",
  1153 => x"87c578c0",
  1154 => x"c148a6cc",
  1155 => x"4966cc78",
  1156 => x"c487ffea",
  1157 => x"6e7e7086",
  1158 => x"87e9c202",
  1159 => x"81cb496e",
  1160 => x"d0496997",
  1161 => x"d6c10299",
  1162 => x"e7c5c187",
  1163 => x"cb49744a",
  1164 => x"d3e8c191",
  1165 => x"c8797281",
  1166 => x"51ffc381",
  1167 => x"91de4974",
  1168 => x"4dd1dec3",
  1169 => x"c1c28571",
  1170 => x"a5c17d97",
  1171 => x"51e0c049",
  1172 => x"97d6d9c3",
  1173 => x"87d202bf",
  1174 => x"a5c284c1",
  1175 => x"d6d9c34b",
  1176 => x"fe49db4a",
  1177 => x"c187c1f9",
  1178 => x"a5cd87db",
  1179 => x"c151c049",
  1180 => x"4ba5c284",
  1181 => x"49cb4a6e",
  1182 => x"87ecf8fe",
  1183 => x"c187c6c1",
  1184 => x"744ae3c3",
  1185 => x"c191cb49",
  1186 => x"7281d3e8",
  1187 => x"d6d9c379",
  1188 => x"d802bf97",
  1189 => x"de497487",
  1190 => x"c384c191",
  1191 => x"714bd1de",
  1192 => x"d6d9c383",
  1193 => x"fe49dd4a",
  1194 => x"d887fdf7",
  1195 => x"de4b7487",
  1196 => x"d1dec393",
  1197 => x"49a3cb83",
  1198 => x"84c151c0",
  1199 => x"cb4a6e73",
  1200 => x"e3f7fe49",
  1201 => x"4866c487",
  1202 => x"a6c880c1",
  1203 => x"03acc758",
  1204 => x"6e87c5c0",
  1205 => x"87e0fc05",
  1206 => x"8ef44874",
  1207 => x"1e87fcf7",
  1208 => x"4b711e73",
  1209 => x"c191cb49",
  1210 => x"c881d3e8",
  1211 => x"ccc34aa1",
  1212 => x"501248d5",
  1213 => x"c14aa1c9",
  1214 => x"1248dec2",
  1215 => x"c381ca50",
  1216 => x"1148d0de",
  1217 => x"d0dec350",
  1218 => x"1e49bf97",
  1219 => x"ffc149c0",
  1220 => x"ddc387cc",
  1221 => x"78de48f8",
  1222 => x"cad649c1",
  1223 => x"fef62687",
  1224 => x"4a711e87",
  1225 => x"c191cb49",
  1226 => x"c881d3e8",
  1227 => x"c3481181",
  1228 => x"c358fcdd",
  1229 => x"c048fcdd",
  1230 => x"d549c178",
  1231 => x"4f2687e9",
  1232 => x"c149c01e",
  1233 => x"2687fec1",
  1234 => x"99711e4f",
  1235 => x"c187d202",
  1236 => x"c048e8e9",
  1237 => x"c180f750",
  1238 => x"c140e1cc",
  1239 => x"ce78cce8",
  1240 => x"e4e9c187",
  1241 => x"c5e8c148",
  1242 => x"c180fc78",
  1243 => x"2678c0cd",
  1244 => x"5b5e0e4f",
  1245 => x"4c710e5c",
  1246 => x"c192cb4a",
  1247 => x"c882d3e8",
  1248 => x"a2c949a2",
  1249 => x"4b6b974b",
  1250 => x"4969971e",
  1251 => x"1282ca1e",
  1252 => x"f7eac049",
  1253 => x"d449c087",
  1254 => x"497487cd",
  1255 => x"87c0ffc0",
  1256 => x"f8f48ef8",
  1257 => x"1e731e87",
  1258 => x"ff494b71",
  1259 => x"497387c3",
  1260 => x"c087fefe",
  1261 => x"ccc0c149",
  1262 => x"87e3f487",
  1263 => x"711e731e",
  1264 => x"4aa3c64b",
  1265 => x"c187db02",
  1266 => x"87d6028a",
  1267 => x"dac1028a",
  1268 => x"c0028a87",
  1269 => x"028a87fc",
  1270 => x"8a87e1c0",
  1271 => x"c187cb02",
  1272 => x"49c787db",
  1273 => x"c187fafc",
  1274 => x"ddc387de",
  1275 => x"c102bffc",
  1276 => x"c14887cb",
  1277 => x"c0dec388",
  1278 => x"87c1c158",
  1279 => x"bfc0dec3",
  1280 => x"87f9c002",
  1281 => x"bffcddc3",
  1282 => x"c380c148",
  1283 => x"c058c0de",
  1284 => x"ddc387eb",
  1285 => x"c649bffc",
  1286 => x"c0dec389",
  1287 => x"a9b7c059",
  1288 => x"c387da03",
  1289 => x"c048fcdd",
  1290 => x"c387d278",
  1291 => x"02bfc0de",
  1292 => x"ddc387cb",
  1293 => x"c648bffc",
  1294 => x"c0dec380",
  1295 => x"d149c058",
  1296 => x"497387e5",
  1297 => x"87d8fcc0",
  1298 => x"0e87d4f2",
  1299 => x"0e5c5b5e",
  1300 => x"66cc4c71",
  1301 => x"cb4b741e",
  1302 => x"d3e8c193",
  1303 => x"4aa3c483",
  1304 => x"f1fe496a",
  1305 => x"cbc187d2",
  1306 => x"a3c87bdf",
  1307 => x"5166d449",
  1308 => x"d849a3c9",
  1309 => x"a3ca5166",
  1310 => x"5166dc49",
  1311 => x"87ddf126",
  1312 => x"5c5b5e0e",
  1313 => x"d0ff0e5d",
  1314 => x"59a6d886",
  1315 => x"c048a6c4",
  1316 => x"c180c478",
  1317 => x"c47866c4",
  1318 => x"c478c180",
  1319 => x"c378c180",
  1320 => x"c148c0de",
  1321 => x"f8ddc378",
  1322 => x"a8de48bf",
  1323 => x"f387cb05",
  1324 => x"497087df",
  1325 => x"ce59a6c8",
  1326 => x"d6e887f6",
  1327 => x"87f8e887",
  1328 => x"7087c5e8",
  1329 => x"acfbc04c",
  1330 => x"87d0c102",
  1331 => x"c10566d4",
  1332 => x"1ec087c2",
  1333 => x"c11ec11e",
  1334 => x"c01ef6e9",
  1335 => x"87ebfd49",
  1336 => x"4a66d0c1",
  1337 => x"496a82c4",
  1338 => x"517481c7",
  1339 => x"1ed81ec1",
  1340 => x"81c8496a",
  1341 => x"d887d5e8",
  1342 => x"66c4c186",
  1343 => x"01a8c048",
  1344 => x"a6c487c7",
  1345 => x"ce78c148",
  1346 => x"66c4c187",
  1347 => x"cc88c148",
  1348 => x"87c358a6",
  1349 => x"cc87e1e7",
  1350 => x"78c248a6",
  1351 => x"cd029c74",
  1352 => x"66c487ca",
  1353 => x"66c8c148",
  1354 => x"ffcc03a8",
  1355 => x"48a6d887",
  1356 => x"d3e678c0",
  1357 => x"c14c7087",
  1358 => x"c205acd0",
  1359 => x"66d887d6",
  1360 => x"87f7e87e",
  1361 => x"a6dc4970",
  1362 => x"87fce559",
  1363 => x"ecc04c70",
  1364 => x"eac105ac",
  1365 => x"4966c487",
  1366 => x"c0c191cb",
  1367 => x"a1c48166",
  1368 => x"c84d6a4a",
  1369 => x"66d84aa1",
  1370 => x"e1ccc152",
  1371 => x"87d8e579",
  1372 => x"029c4c70",
  1373 => x"fbc087d8",
  1374 => x"87d202ac",
  1375 => x"c7e55574",
  1376 => x"9c4c7087",
  1377 => x"c087c702",
  1378 => x"ff05acfb",
  1379 => x"e0c087ee",
  1380 => x"55c1c255",
  1381 => x"d47d97c0",
  1382 => x"a96e4966",
  1383 => x"c487db05",
  1384 => x"66c84866",
  1385 => x"87ca04a8",
  1386 => x"c14866c4",
  1387 => x"58a6c880",
  1388 => x"66c887c8",
  1389 => x"cc88c148",
  1390 => x"cbe458a6",
  1391 => x"c14c7087",
  1392 => x"c805acd0",
  1393 => x"4866d087",
  1394 => x"a6d480c1",
  1395 => x"acd0c158",
  1396 => x"87eafd02",
  1397 => x"d448a6dc",
  1398 => x"66d87866",
  1399 => x"a866dc48",
  1400 => x"87dac905",
  1401 => x"48a6e0c0",
  1402 => x"c478f0c0",
  1403 => x"7866cc80",
  1404 => x"78c080c4",
  1405 => x"c048747e",
  1406 => x"f0c088fb",
  1407 => x"987058a6",
  1408 => x"87d5c802",
  1409 => x"c088cb48",
  1410 => x"7058a6f0",
  1411 => x"e9c00298",
  1412 => x"88c94887",
  1413 => x"58a6f0c0",
  1414 => x"c3029870",
  1415 => x"c44887e1",
  1416 => x"a6f0c088",
  1417 => x"02987058",
  1418 => x"c14887d6",
  1419 => x"a6f0c088",
  1420 => x"02987058",
  1421 => x"c787c8c3",
  1422 => x"e0c087d9",
  1423 => x"78c048a6",
  1424 => x"c14866cc",
  1425 => x"58a6d080",
  1426 => x"7087fde1",
  1427 => x"acecc04c",
  1428 => x"c087d502",
  1429 => x"c60266e0",
  1430 => x"a6e4c087",
  1431 => x"7487c95c",
  1432 => x"88f0c048",
  1433 => x"58a6e8c0",
  1434 => x"02acecc0",
  1435 => x"d7e187cc",
  1436 => x"c04c7087",
  1437 => x"ff05acec",
  1438 => x"e0c087f4",
  1439 => x"66d41e66",
  1440 => x"ecc01e49",
  1441 => x"e9c11e66",
  1442 => x"66d41ef6",
  1443 => x"87fbf649",
  1444 => x"1eca1ec0",
  1445 => x"cb4966dc",
  1446 => x"66d8c191",
  1447 => x"48a6d881",
  1448 => x"d878a1c4",
  1449 => x"e149bf66",
  1450 => x"86d887e2",
  1451 => x"06a8b7c0",
  1452 => x"c187c7c1",
  1453 => x"c81ede1e",
  1454 => x"e149bf66",
  1455 => x"86c887ce",
  1456 => x"c0484970",
  1457 => x"e4c08808",
  1458 => x"b7c058a6",
  1459 => x"e9c006a8",
  1460 => x"66e0c087",
  1461 => x"a8b7dd48",
  1462 => x"6e87df03",
  1463 => x"e0c049bf",
  1464 => x"e0c08166",
  1465 => x"c1496651",
  1466 => x"81bf6e81",
  1467 => x"c051c1c2",
  1468 => x"c24966e0",
  1469 => x"81bf6e81",
  1470 => x"7ec151c0",
  1471 => x"e187dac4",
  1472 => x"e4c087f9",
  1473 => x"f2e158a6",
  1474 => x"a6e8c087",
  1475 => x"a8ecc058",
  1476 => x"87cbc005",
  1477 => x"48a6e4c0",
  1478 => x"7866e0c0",
  1479 => x"ff87c4c0",
  1480 => x"c487e5de",
  1481 => x"91cb4966",
  1482 => x"4866c0c1",
  1483 => x"7e708071",
  1484 => x"81c8496e",
  1485 => x"82ca4a6e",
  1486 => x"5266e0c0",
  1487 => x"4a66e4c0",
  1488 => x"e0c082c1",
  1489 => x"48c18a66",
  1490 => x"4a703072",
  1491 => x"97728ac1",
  1492 => x"49699779",
  1493 => x"66e4c01e",
  1494 => x"87f2da49",
  1495 => x"f0c086c4",
  1496 => x"496e58a6",
  1497 => x"4d6981c4",
  1498 => x"d84866dc",
  1499 => x"c002a866",
  1500 => x"a6d887c8",
  1501 => x"c078c048",
  1502 => x"a6d887c5",
  1503 => x"d878c148",
  1504 => x"e0c01e66",
  1505 => x"ff49751e",
  1506 => x"c887c1de",
  1507 => x"c04c7086",
  1508 => x"c106acb7",
  1509 => x"857487d4",
  1510 => x"7449e0c0",
  1511 => x"c14b7589",
  1512 => x"714ae4e2",
  1513 => x"87c0e4fe",
  1514 => x"e8c085c2",
  1515 => x"80c14866",
  1516 => x"58a6ecc0",
  1517 => x"4966ecc0",
  1518 => x"a97081c1",
  1519 => x"87c8c002",
  1520 => x"c048a6d8",
  1521 => x"87c5c078",
  1522 => x"c148a6d8",
  1523 => x"1e66d878",
  1524 => x"c049a4c2",
  1525 => x"887148e0",
  1526 => x"751e4970",
  1527 => x"ebdcff49",
  1528 => x"c086c887",
  1529 => x"ff01a8b7",
  1530 => x"e8c087c0",
  1531 => x"d1c00266",
  1532 => x"c9496e87",
  1533 => x"66e8c081",
  1534 => x"c1486e51",
  1535 => x"c078f1cd",
  1536 => x"496e87cc",
  1537 => x"51c281c9",
  1538 => x"cec1486e",
  1539 => x"7ec178e5",
  1540 => x"ff87c6c0",
  1541 => x"7087e1db",
  1542 => x"c0026e4c",
  1543 => x"66c487f5",
  1544 => x"a866c848",
  1545 => x"87cbc004",
  1546 => x"c14866c4",
  1547 => x"58a6c880",
  1548 => x"c887e0c0",
  1549 => x"88c14866",
  1550 => x"c058a6cc",
  1551 => x"c6c187d5",
  1552 => x"c8c005ac",
  1553 => x"4866cc87",
  1554 => x"a6d080c1",
  1555 => x"e7daff58",
  1556 => x"d04c7087",
  1557 => x"80c14866",
  1558 => x"7458a6d4",
  1559 => x"cbc0029c",
  1560 => x"4866c487",
  1561 => x"a866c8c1",
  1562 => x"87c1f304",
  1563 => x"87ffd9ff",
  1564 => x"c74866c4",
  1565 => x"e5c003a8",
  1566 => x"c0dec387",
  1567 => x"c478c048",
  1568 => x"91cb4966",
  1569 => x"8166c0c1",
  1570 => x"6a4aa1c4",
  1571 => x"7952c04a",
  1572 => x"c14866c4",
  1573 => x"58a6c880",
  1574 => x"ff04a8c7",
  1575 => x"d0ff87db",
  1576 => x"87f7e08e",
  1577 => x"1e00203a",
  1578 => x"4b711e73",
  1579 => x"87c6029b",
  1580 => x"48fcddc3",
  1581 => x"1ec778c0",
  1582 => x"bffcddc3",
  1583 => x"e8c11e49",
  1584 => x"ddc31ed3",
  1585 => x"ee49bff8",
  1586 => x"86cc87f6",
  1587 => x"bff8ddc3",
  1588 => x"87f5e949",
  1589 => x"c8029b73",
  1590 => x"d3e8c187",
  1591 => x"d1ebc049",
  1592 => x"fadfff87",
  1593 => x"1e731e87",
  1594 => x"4bffc31e",
  1595 => x"fc4ad4ff",
  1596 => x"98c148bf",
  1597 => x"026e7e70",
  1598 => x"ff87fbc0",
  1599 => x"c1c148d0",
  1600 => x"7ad2c278",
  1601 => x"d1c37a73",
  1602 => x"ff4849c7",
  1603 => x"73506a80",
  1604 => x"73516a7a",
  1605 => x"6a80c17a",
  1606 => x"6a7a7350",
  1607 => x"6a7a7350",
  1608 => x"6a7a7349",
  1609 => x"6a7a7350",
  1610 => x"d0d1c350",
  1611 => x"d0ff5997",
  1612 => x"78c0c148",
  1613 => x"d1c387d7",
  1614 => x"ff4849c7",
  1615 => x"5150c080",
  1616 => x"50c080c1",
  1617 => x"50c150d9",
  1618 => x"c350e2c0",
  1619 => x"cdd1c350",
  1620 => x"f850c048",
  1621 => x"deff2680",
  1622 => x"c71e87c5",
  1623 => x"49c187f7",
  1624 => x"fe87c4fd",
  1625 => x"7087c6e7",
  1626 => x"87cd0298",
  1627 => x"87c3f0fe",
  1628 => x"c4029870",
  1629 => x"c24ac187",
  1630 => x"724ac087",
  1631 => x"87ce059a",
  1632 => x"e6c11ec0",
  1633 => x"f5c049ef",
  1634 => x"86c487f7",
  1635 => x"e6c187fe",
  1636 => x"1ec087ed",
  1637 => x"49fae6c1",
  1638 => x"87e5f5c0",
  1639 => x"e7c11ec0",
  1640 => x"497087c6",
  1641 => x"87d9f5c0",
  1642 => x"f887e9c3",
  1643 => x"534f268e",
  1644 => x"61662044",
  1645 => x"64656c69",
  1646 => x"6f42002e",
  1647 => x"6e69746f",
  1648 => x"2e2e2e67",
  1649 => x"c01e1e00",
  1650 => x"c187c3ec",
  1651 => x"6e87dcda",
  1652 => x"ffffc149",
  1653 => x"c1486e99",
  1654 => x"717e7080",
  1655 => x"87e70599",
  1656 => x"7087c2fc",
  1657 => x"87f5ce49",
  1658 => x"2687dcff",
  1659 => x"c31e4f26",
  1660 => x"c048fcdd",
  1661 => x"f8ddc378",
  1662 => x"fd78c048",
  1663 => x"c4ff87dc",
  1664 => x"2648c087",
  1665 => x"4520804f",
  1666 => x"00746978",
  1667 => x"61422080",
  1668 => x"21006b63",
  1669 => x"91000013",
  1670 => x"00000037",
  1671 => x"13210000",
  1672 => x"37af0000",
  1673 => x"00000000",
  1674 => x"00132100",
  1675 => x"0037cd00",
  1676 => x"00000000",
  1677 => x"00001321",
  1678 => x"000037eb",
  1679 => x"21000000",
  1680 => x"09000013",
  1681 => x"00000038",
  1682 => x"13210000",
  1683 => x"38270000",
  1684 => x"00000000",
  1685 => x"00132100",
  1686 => x"00384500",
  1687 => x"00000000",
  1688 => x"00001321",
  1689 => x"00000000",
  1690 => x"bc000000",
  1691 => x"00000013",
  1692 => x"00000000",
  1693 => x"6f4c0000",
  1694 => x"2a206461",
  1695 => x"fe1e002e",
  1696 => x"78c048f0",
  1697 => x"097909cd",
  1698 => x"1e1e4f26",
  1699 => x"7ebff0fe",
  1700 => x"4f262648",
  1701 => x"48f0fe1e",
  1702 => x"4f2678c1",
  1703 => x"48f0fe1e",
  1704 => x"4f2678c0",
  1705 => x"c04a711e",
  1706 => x"4f265252",
  1707 => x"5c5b5e0e",
  1708 => x"86f40e5d",
  1709 => x"6d974d71",
  1710 => x"4ca5c17e",
  1711 => x"c8486c97",
  1712 => x"486e58a6",
  1713 => x"05a866c4",
  1714 => x"48ff87c5",
  1715 => x"ff87e6c0",
  1716 => x"a5c287ca",
  1717 => x"4b6c9749",
  1718 => x"974ba371",
  1719 => x"6c974b6b",
  1720 => x"c1486e7e",
  1721 => x"58a6c880",
  1722 => x"a6cc98c7",
  1723 => x"7c977058",
  1724 => x"7387e1fe",
  1725 => x"268ef448",
  1726 => x"264c264d",
  1727 => x"0e4f264b",
  1728 => x"0e5c5b5e",
  1729 => x"4c7186f4",
  1730 => x"c34a66d8",
  1731 => x"a4c29aff",
  1732 => x"496c974b",
  1733 => x"7249a173",
  1734 => x"7e6c9751",
  1735 => x"80c1486e",
  1736 => x"c758a6c8",
  1737 => x"58a6cc98",
  1738 => x"8ef45470",
  1739 => x"1e87caff",
  1740 => x"87e8fd1e",
  1741 => x"494abfe0",
  1742 => x"99c0e0c0",
  1743 => x"7287cb02",
  1744 => x"e3e1c31e",
  1745 => x"87f7fe49",
  1746 => x"fdfc86c4",
  1747 => x"fd7e7087",
  1748 => x"262687c2",
  1749 => x"e1c31e4f",
  1750 => x"c7fd49e3",
  1751 => x"efecc187",
  1752 => x"87dafc49",
  1753 => x"2687d9c5",
  1754 => x"5b5e0e4f",
  1755 => x"c30e5d5c",
  1756 => x"4abfc6e2",
  1757 => x"bffdeec1",
  1758 => x"bc724c49",
  1759 => x"dbfc4d71",
  1760 => x"744bc087",
  1761 => x"0299d049",
  1762 => x"497587d5",
  1763 => x"1e7199d0",
  1764 => x"f5c11ec0",
  1765 => x"82734acf",
  1766 => x"e4c04912",
  1767 => x"c186c887",
  1768 => x"c8832d2c",
  1769 => x"daff04ab",
  1770 => x"87e8fb87",
  1771 => x"48fdeec1",
  1772 => x"bfc6e2c3",
  1773 => x"264d2678",
  1774 => x"264b264c",
  1775 => x"0000004f",
  1776 => x"d0ff1e00",
  1777 => x"78e1c848",
  1778 => x"c548d4ff",
  1779 => x"0266c478",
  1780 => x"e0c387c3",
  1781 => x"0266c878",
  1782 => x"d4ff87c6",
  1783 => x"78f0c348",
  1784 => x"7148d4ff",
  1785 => x"48d0ff78",
  1786 => x"c078e1c8",
  1787 => x"4f2678e0",
  1788 => x"5c5b5e0e",
  1789 => x"c34c710e",
  1790 => x"fa49e3e1",
  1791 => x"4a7087ee",
  1792 => x"04aab7c0",
  1793 => x"c387e3c2",
  1794 => x"c905aae0",
  1795 => x"f3f2c187",
  1796 => x"c278c148",
  1797 => x"f0c387d4",
  1798 => x"87c905aa",
  1799 => x"48eff2c1",
  1800 => x"f5c178c1",
  1801 => x"f3f2c187",
  1802 => x"87c702bf",
  1803 => x"c0c24b72",
  1804 => x"7287c2b3",
  1805 => x"059c744b",
  1806 => x"f2c187d1",
  1807 => x"c11ebfef",
  1808 => x"1ebff3f2",
  1809 => x"f8fd4972",
  1810 => x"c186c887",
  1811 => x"02bfeff2",
  1812 => x"7387e0c0",
  1813 => x"29b7c449",
  1814 => x"cff4c191",
  1815 => x"cf4a7381",
  1816 => x"c192c29a",
  1817 => x"70307248",
  1818 => x"72baff4a",
  1819 => x"70986948",
  1820 => x"7387db79",
  1821 => x"29b7c449",
  1822 => x"cff4c191",
  1823 => x"cf4a7381",
  1824 => x"c392c29a",
  1825 => x"70307248",
  1826 => x"b069484a",
  1827 => x"f2c17970",
  1828 => x"78c048f3",
  1829 => x"48eff2c1",
  1830 => x"e1c378c0",
  1831 => x"cbf849e3",
  1832 => x"c04a7087",
  1833 => x"fd03aab7",
  1834 => x"48c087dd",
  1835 => x"0087c8fc",
  1836 => x"00000000",
  1837 => x"1e000000",
  1838 => x"fc494a71",
  1839 => x"4f2687f2",
  1840 => x"724ac01e",
  1841 => x"c191c449",
  1842 => x"c081cff4",
  1843 => x"d082c179",
  1844 => x"ee04aab7",
  1845 => x"0e4f2687",
  1846 => x"5d5c5b5e",
  1847 => x"f64d710e",
  1848 => x"4a7587fa",
  1849 => x"922ab7c4",
  1850 => x"82cff4c1",
  1851 => x"9ccf4c75",
  1852 => x"496a94c2",
  1853 => x"c32b744b",
  1854 => x"7448c29b",
  1855 => x"ff4c7030",
  1856 => x"714874bc",
  1857 => x"f67a7098",
  1858 => x"487387ca",
  1859 => x"0087e6fa",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"00000000",
  1868 => x"00000000",
  1869 => x"00000000",
  1870 => x"00000000",
  1871 => x"00000000",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00000000",
  1875 => x"16000000",
  1876 => x"2e25261e",
  1877 => x"1e3e3d36",
  1878 => x"c848d0ff",
  1879 => x"487178e1",
  1880 => x"7808d4ff",
  1881 => x"ff1e4f26",
  1882 => x"e1c848d0",
  1883 => x"ff487178",
  1884 => x"c47808d4",
  1885 => x"d4ff4866",
  1886 => x"4f267808",
  1887 => x"c44a711e",
  1888 => x"e0c11e66",
  1889 => x"ddff49a2",
  1890 => x"4966c887",
  1891 => x"ff29b7c8",
  1892 => x"787148d4",
  1893 => x"c048d0ff",
  1894 => x"262678e0",
  1895 => x"1e731e4f",
  1896 => x"e2c04b71",
  1897 => x"87effe49",
  1898 => x"48134ac7",
  1899 => x"7808d4ff",
  1900 => x"8ac14972",
  1901 => x"f1059971",
  1902 => x"48d0ff87",
  1903 => x"c478e0c0",
  1904 => x"264d2687",
  1905 => x"264b264c",
  1906 => x"d4ff1e4f",
  1907 => x"7affc34a",
  1908 => x"c848d0ff",
  1909 => x"7ade78e1",
  1910 => x"bfede1c3",
  1911 => x"c848497a",
  1912 => x"717a7028",
  1913 => x"7028d048",
  1914 => x"d848717a",
  1915 => x"c37a7028",
  1916 => x"7abff1e1",
  1917 => x"28c84849",
  1918 => x"48717a70",
  1919 => x"7a7028d0",
  1920 => x"28d84871",
  1921 => x"d0ff7a70",
  1922 => x"78e0c048",
  1923 => x"731e4f26",
  1924 => x"c34a711e",
  1925 => x"4bbfede1",
  1926 => x"e0c02b72",
  1927 => x"87ce04aa",
  1928 => x"e0c04972",
  1929 => x"f1e1c389",
  1930 => x"2b714bbf",
  1931 => x"e0c087cf",
  1932 => x"c3897249",
  1933 => x"48bff1e1",
  1934 => x"49703071",
  1935 => x"9b66c8b3",
  1936 => x"87c44873",
  1937 => x"4c264d26",
  1938 => x"4f264b26",
  1939 => x"5c5b5e0e",
  1940 => x"86ec0e5d",
  1941 => x"e1c34b71",
  1942 => x"4c7ebfed",
  1943 => x"e0c02c73",
  1944 => x"e0c004ab",
  1945 => x"48a6c487",
  1946 => x"497378c0",
  1947 => x"7189e0c0",
  1948 => x"66e4c04a",
  1949 => x"cc307248",
  1950 => x"e1c358a6",
  1951 => x"4c4dbff1",
  1952 => x"e4c02c71",
  1953 => x"c0497387",
  1954 => x"714866e4",
  1955 => x"58a6c830",
  1956 => x"7349e0c0",
  1957 => x"66e4c089",
  1958 => x"cc287148",
  1959 => x"e1c358a6",
  1960 => x"484dbff1",
  1961 => x"49703071",
  1962 => x"66e4c0b4",
  1963 => x"c084c19c",
  1964 => x"04ac66e8",
  1965 => x"4cc087c2",
  1966 => x"04abe0c0",
  1967 => x"a6cc87d3",
  1968 => x"7378c048",
  1969 => x"89e0c049",
  1970 => x"30714874",
  1971 => x"d558a6d4",
  1972 => x"74497387",
  1973 => x"d0307148",
  1974 => x"e0c058a6",
  1975 => x"74897349",
  1976 => x"d4287148",
  1977 => x"66c458a6",
  1978 => x"6ebaff4a",
  1979 => x"4966c89a",
  1980 => x"9975b9ff",
  1981 => x"66cc4872",
  1982 => x"f1e1c3b0",
  1983 => x"d0487158",
  1984 => x"e1c3b066",
  1985 => x"c0fb58f5",
  1986 => x"fc8eec87",
  1987 => x"ff1e87f6",
  1988 => x"c9c848d0",
  1989 => x"ff487178",
  1990 => x"267808d4",
  1991 => x"4a711e4f",
  1992 => x"ff87eb49",
  1993 => x"78c848d0",
  1994 => x"731e4f26",
  1995 => x"c34b711e",
  1996 => x"02bfc1e2",
  1997 => x"ebc287c3",
  1998 => x"48d0ff87",
  1999 => x"7378c9c8",
  2000 => x"b1e0c049",
  2001 => x"7148d4ff",
  2002 => x"f5e1c378",
  2003 => x"c878c048",
  2004 => x"87c50266",
  2005 => x"c249ffc3",
  2006 => x"c349c087",
  2007 => x"cc59fde1",
  2008 => x"87c60266",
  2009 => x"4ad5d5c5",
  2010 => x"ffcf87c4",
  2011 => x"e2c34aff",
  2012 => x"e2c35ac1",
  2013 => x"78c148c1",
  2014 => x"4d2687c4",
  2015 => x"4b264c26",
  2016 => x"5e0e4f26",
  2017 => x"0e5d5c5b",
  2018 => x"e1c34a71",
  2019 => x"724cbffd",
  2020 => x"87cb029a",
  2021 => x"c191c849",
  2022 => x"714be0fc",
  2023 => x"c287c483",
  2024 => x"c04be0c0",
  2025 => x"7449134d",
  2026 => x"f9e1c399",
  2027 => x"d4ffb9bf",
  2028 => x"c1787148",
  2029 => x"c8852cb7",
  2030 => x"e804adb7",
  2031 => x"f5e1c387",
  2032 => x"80c848bf",
  2033 => x"58f9e1c3",
  2034 => x"1e87effe",
  2035 => x"4b711e73",
  2036 => x"029a4a13",
  2037 => x"497287cb",
  2038 => x"1387e7fe",
  2039 => x"f5059a4a",
  2040 => x"87dafe87",
  2041 => x"f5e1c31e",
  2042 => x"e1c349bf",
  2043 => x"a1c148f5",
  2044 => x"b7c0c478",
  2045 => x"87db03a9",
  2046 => x"c348d4ff",
  2047 => x"78bff9e1",
  2048 => x"bff5e1c3",
  2049 => x"f5e1c349",
  2050 => x"78a1c148",
  2051 => x"a9b7c0c4",
  2052 => x"ff87e504",
  2053 => x"78c848d0",
  2054 => x"48c1e2c3",
  2055 => x"4f2678c0",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"5f000000",
  2059 => x"0000005f",
  2060 => x"00030300",
  2061 => x"00000303",
  2062 => x"147f7f14",
  2063 => x"00147f7f",
  2064 => x"6b2e2400",
  2065 => x"00123a6b",
  2066 => x"18366a4c",
  2067 => x"0032566c",
  2068 => x"594f7e30",
  2069 => x"40683a77",
  2070 => x"07040000",
  2071 => x"00000003",
  2072 => x"3e1c0000",
  2073 => x"00004163",
  2074 => x"63410000",
  2075 => x"00001c3e",
  2076 => x"1c3e2a08",
  2077 => x"082a3e1c",
  2078 => x"3e080800",
  2079 => x"0008083e",
  2080 => x"e0800000",
  2081 => x"00000060",
  2082 => x"08080800",
  2083 => x"00080808",
  2084 => x"60000000",
  2085 => x"00000060",
  2086 => x"18306040",
  2087 => x"0103060c",
  2088 => x"597f3e00",
  2089 => x"003e7f4d",
  2090 => x"7f060400",
  2091 => x"0000007f",
  2092 => x"71634200",
  2093 => x"00464f59",
  2094 => x"49632200",
  2095 => x"00367f49",
  2096 => x"13161c18",
  2097 => x"00107f7f",
  2098 => x"45672700",
  2099 => x"00397d45",
  2100 => x"4b7e3c00",
  2101 => x"00307949",
  2102 => x"71010100",
  2103 => x"00070f79",
  2104 => x"497f3600",
  2105 => x"00367f49",
  2106 => x"494f0600",
  2107 => x"001e3f69",
  2108 => x"66000000",
  2109 => x"00000066",
  2110 => x"e6800000",
  2111 => x"00000066",
  2112 => x"14080800",
  2113 => x"00222214",
  2114 => x"14141400",
  2115 => x"00141414",
  2116 => x"14222200",
  2117 => x"00080814",
  2118 => x"51030200",
  2119 => x"00060f59",
  2120 => x"5d417f3e",
  2121 => x"001e1f55",
  2122 => x"097f7e00",
  2123 => x"007e7f09",
  2124 => x"497f7f00",
  2125 => x"00367f49",
  2126 => x"633e1c00",
  2127 => x"00414141",
  2128 => x"417f7f00",
  2129 => x"001c3e63",
  2130 => x"497f7f00",
  2131 => x"00414149",
  2132 => x"097f7f00",
  2133 => x"00010109",
  2134 => x"417f3e00",
  2135 => x"007a7b49",
  2136 => x"087f7f00",
  2137 => x"007f7f08",
  2138 => x"7f410000",
  2139 => x"0000417f",
  2140 => x"40602000",
  2141 => x"003f7f40",
  2142 => x"1c087f7f",
  2143 => x"00416336",
  2144 => x"407f7f00",
  2145 => x"00404040",
  2146 => x"0c067f7f",
  2147 => x"007f7f06",
  2148 => x"0c067f7f",
  2149 => x"007f7f18",
  2150 => x"417f3e00",
  2151 => x"003e7f41",
  2152 => x"097f7f00",
  2153 => x"00060f09",
  2154 => x"61417f3e",
  2155 => x"00407e7f",
  2156 => x"097f7f00",
  2157 => x"00667f19",
  2158 => x"4d6f2600",
  2159 => x"00327b59",
  2160 => x"7f010100",
  2161 => x"0001017f",
  2162 => x"407f3f00",
  2163 => x"003f7f40",
  2164 => x"703f0f00",
  2165 => x"000f3f70",
  2166 => x"18307f7f",
  2167 => x"007f7f30",
  2168 => x"1c366341",
  2169 => x"4163361c",
  2170 => x"7c060301",
  2171 => x"0103067c",
  2172 => x"4d597161",
  2173 => x"00414347",
  2174 => x"7f7f0000",
  2175 => x"00004141",
  2176 => x"0c060301",
  2177 => x"40603018",
  2178 => x"41410000",
  2179 => x"00007f7f",
  2180 => x"03060c08",
  2181 => x"00080c06",
  2182 => x"80808080",
  2183 => x"00808080",
  2184 => x"03000000",
  2185 => x"00000407",
  2186 => x"54742000",
  2187 => x"00787c54",
  2188 => x"447f7f00",
  2189 => x"00387c44",
  2190 => x"447c3800",
  2191 => x"00004444",
  2192 => x"447c3800",
  2193 => x"007f7f44",
  2194 => x"547c3800",
  2195 => x"00185c54",
  2196 => x"7f7e0400",
  2197 => x"00000505",
  2198 => x"a4bc1800",
  2199 => x"007cfca4",
  2200 => x"047f7f00",
  2201 => x"00787c04",
  2202 => x"3d000000",
  2203 => x"0000407d",
  2204 => x"80808000",
  2205 => x"00007dfd",
  2206 => x"107f7f00",
  2207 => x"00446c38",
  2208 => x"3f000000",
  2209 => x"0000407f",
  2210 => x"180c7c7c",
  2211 => x"00787c0c",
  2212 => x"047c7c00",
  2213 => x"00787c04",
  2214 => x"447c3800",
  2215 => x"00387c44",
  2216 => x"24fcfc00",
  2217 => x"00183c24",
  2218 => x"243c1800",
  2219 => x"00fcfc24",
  2220 => x"047c7c00",
  2221 => x"00080c04",
  2222 => x"545c4800",
  2223 => x"00207454",
  2224 => x"7f3f0400",
  2225 => x"00004444",
  2226 => x"407c3c00",
  2227 => x"007c7c40",
  2228 => x"603c1c00",
  2229 => x"001c3c60",
  2230 => x"30607c3c",
  2231 => x"003c7c60",
  2232 => x"10386c44",
  2233 => x"00446c38",
  2234 => x"e0bc1c00",
  2235 => x"001c3c60",
  2236 => x"74644400",
  2237 => x"00444c5c",
  2238 => x"3e080800",
  2239 => x"00414177",
  2240 => x"7f000000",
  2241 => x"0000007f",
  2242 => x"77414100",
  2243 => x"0008083e",
  2244 => x"03010102",
  2245 => x"00010202",
  2246 => x"7f7f7f7f",
  2247 => x"007f7f7f",
  2248 => x"1c1c0808",
  2249 => x"7f7f3e3e",
  2250 => x"3e3e7f7f",
  2251 => x"08081c1c",
  2252 => x"7c181000",
  2253 => x"0010187c",
  2254 => x"7c301000",
  2255 => x"0010307c",
  2256 => x"60603010",
  2257 => x"00061e78",
  2258 => x"183c6642",
  2259 => x"0042663c",
  2260 => x"c26a3878",
  2261 => x"00386cc6",
  2262 => x"60000060",
  2263 => x"00600000",
  2264 => x"5c5b5e0e",
  2265 => x"711e0e5d",
  2266 => x"d2e2c34c",
  2267 => x"4bc04dbf",
  2268 => x"ab741ec0",
  2269 => x"c487c702",
  2270 => x"78c048a6",
  2271 => x"a6c487c5",
  2272 => x"c478c148",
  2273 => x"49731e66",
  2274 => x"c887dfee",
  2275 => x"49e0c086",
  2276 => x"c487efef",
  2277 => x"496a4aa5",
  2278 => x"f187f0f0",
  2279 => x"85cb87c6",
  2280 => x"b7c883c1",
  2281 => x"c7ff04ab",
  2282 => x"4d262687",
  2283 => x"4b264c26",
  2284 => x"711e4f26",
  2285 => x"d6e2c34a",
  2286 => x"d6e2c35a",
  2287 => x"4978c748",
  2288 => x"2687ddfe",
  2289 => x"1e731e4f",
  2290 => x"b7c04a71",
  2291 => x"87d303aa",
  2292 => x"bfe7ddc2",
  2293 => x"c187c405",
  2294 => x"c087c24b",
  2295 => x"ebddc24b",
  2296 => x"c287c45b",
  2297 => x"c25aebdd",
  2298 => x"4abfe7dd",
  2299 => x"c0c19ac1",
  2300 => x"e8ec49a2",
  2301 => x"c248fc87",
  2302 => x"78bfe7dd",
  2303 => x"1e87effe",
  2304 => x"66c44a71",
  2305 => x"e549721e",
  2306 => x"262687f2",
  2307 => x"ddc21e4f",
  2308 => x"e249bfe7",
  2309 => x"e2c387e1",
  2310 => x"bfe848ca",
  2311 => x"c6e2c378",
  2312 => x"78bfec48",
  2313 => x"bfcae2c3",
  2314 => x"ffc3494a",
  2315 => x"2ab7c899",
  2316 => x"b0714872",
  2317 => x"58d2e2c3",
  2318 => x"5e0e4f26",
  2319 => x"0e5d5c5b",
  2320 => x"c8ff4b71",
  2321 => x"c5e2c387",
  2322 => x"7350c048",
  2323 => x"87c7e249",
  2324 => x"c24c4970",
  2325 => x"49eecb9c",
  2326 => x"7087d4cc",
  2327 => x"e2c34d49",
  2328 => x"05bf97c5",
  2329 => x"d087e2c1",
  2330 => x"e2c34966",
  2331 => x"0599bfce",
  2332 => x"66d487d6",
  2333 => x"c6e2c349",
  2334 => x"cb0599bf",
  2335 => x"e1497387",
  2336 => x"987087d5",
  2337 => x"87c1c102",
  2338 => x"c0fe4cc1",
  2339 => x"cb497587",
  2340 => x"987087e9",
  2341 => x"c387c602",
  2342 => x"c148c5e2",
  2343 => x"c5e2c350",
  2344 => x"c005bf97",
  2345 => x"e2c387e3",
  2346 => x"d049bfce",
  2347 => x"ff059966",
  2348 => x"e2c387d6",
  2349 => x"d449bfc6",
  2350 => x"ff059966",
  2351 => x"497387ca",
  2352 => x"7087d4e0",
  2353 => x"fffe0598",
  2354 => x"fb487487",
  2355 => x"5e0e87dc",
  2356 => x"0e5d5c5b",
  2357 => x"4dc086f4",
  2358 => x"7ebfec4c",
  2359 => x"c348a6c4",
  2360 => x"78bfd2e2",
  2361 => x"1ec01ec1",
  2362 => x"cdfd49c7",
  2363 => x"7086c887",
  2364 => x"87ce0298",
  2365 => x"ccfb49ff",
  2366 => x"49dac187",
  2367 => x"87d7dfff",
  2368 => x"e2c34dc1",
  2369 => x"02bf97c5",
  2370 => x"f8c087c4",
  2371 => x"e2c387c8",
  2372 => x"c24bbfca",
  2373 => x"05bfe7dd",
  2374 => x"c487dcc1",
  2375 => x"c0c848a6",
  2376 => x"ddc278c0",
  2377 => x"976e7ed3",
  2378 => x"486e49bf",
  2379 => x"7e7080c1",
  2380 => x"e2deff71",
  2381 => x"02987087",
  2382 => x"66c487c3",
  2383 => x"4866c4b3",
  2384 => x"c828b7c1",
  2385 => x"987058a6",
  2386 => x"87daff05",
  2387 => x"ff49fdc3",
  2388 => x"c387c4de",
  2389 => x"ddff49fa",
  2390 => x"497387fd",
  2391 => x"7199ffc3",
  2392 => x"fa49c01e",
  2393 => x"497387d9",
  2394 => x"7129b7c8",
  2395 => x"fa49c11e",
  2396 => x"86c887cd",
  2397 => x"c387c5c6",
  2398 => x"4bbfcee2",
  2399 => x"87dd029b",
  2400 => x"bfe3ddc2",
  2401 => x"87f3c749",
  2402 => x"c4059870",
  2403 => x"d24bc087",
  2404 => x"49e0c287",
  2405 => x"c287d8c7",
  2406 => x"c658e7dd",
  2407 => x"e3ddc287",
  2408 => x"7378c048",
  2409 => x"0599c249",
  2410 => x"ebc387cf",
  2411 => x"e6dcff49",
  2412 => x"c2497087",
  2413 => x"c2c00299",
  2414 => x"734cfb87",
  2415 => x"0599c149",
  2416 => x"f4c387cf",
  2417 => x"cedcff49",
  2418 => x"c2497087",
  2419 => x"c2c00299",
  2420 => x"734cfa87",
  2421 => x"0599c849",
  2422 => x"f5c387ce",
  2423 => x"f6dbff49",
  2424 => x"c2497087",
  2425 => x"87d60299",
  2426 => x"bfd6e2c3",
  2427 => x"87cac002",
  2428 => x"c388c148",
  2429 => x"c058dae2",
  2430 => x"4cff87c2",
  2431 => x"49734dc1",
  2432 => x"c00599c4",
  2433 => x"f2c387ce",
  2434 => x"cadbff49",
  2435 => x"c2497087",
  2436 => x"87dc0299",
  2437 => x"bfd6e2c3",
  2438 => x"b7c7487e",
  2439 => x"cbc003a8",
  2440 => x"c1486e87",
  2441 => x"dae2c380",
  2442 => x"87c2c058",
  2443 => x"4dc14cfe",
  2444 => x"ff49fdc3",
  2445 => x"7087e0da",
  2446 => x"0299c249",
  2447 => x"c387d5c0",
  2448 => x"02bfd6e2",
  2449 => x"c387c9c0",
  2450 => x"c048d6e2",
  2451 => x"87c2c078",
  2452 => x"4dc14cfd",
  2453 => x"ff49fac3",
  2454 => x"7087fcd9",
  2455 => x"0299c249",
  2456 => x"c387d9c0",
  2457 => x"48bfd6e2",
  2458 => x"03a8b7c7",
  2459 => x"c387c9c0",
  2460 => x"c748d6e2",
  2461 => x"87c2c078",
  2462 => x"4dc14cfc",
  2463 => x"03acb7c0",
  2464 => x"c487d1c0",
  2465 => x"d8c14a66",
  2466 => x"c0026a82",
  2467 => x"4b6a87c6",
  2468 => x"0f734974",
  2469 => x"f0c31ec0",
  2470 => x"49dac11e",
  2471 => x"c887dbf6",
  2472 => x"02987086",
  2473 => x"c887e2c0",
  2474 => x"e2c348a6",
  2475 => x"c878bfd6",
  2476 => x"91cb4966",
  2477 => x"714866c4",
  2478 => x"6e7e7080",
  2479 => x"c8c002bf",
  2480 => x"4bbf6e87",
  2481 => x"734966c8",
  2482 => x"029d750f",
  2483 => x"c387c8c0",
  2484 => x"49bfd6e2",
  2485 => x"c287c9f2",
  2486 => x"02bfebdd",
  2487 => x"4987ddc0",
  2488 => x"7087d8c2",
  2489 => x"d3c00298",
  2490 => x"d6e2c387",
  2491 => x"eff149bf",
  2492 => x"f349c087",
  2493 => x"ddc287cf",
  2494 => x"78c048eb",
  2495 => x"e9f28ef4",
  2496 => x"5b5e0e87",
  2497 => x"1e0e5d5c",
  2498 => x"e2c34c71",
  2499 => x"c149bfd2",
  2500 => x"c14da1cd",
  2501 => x"7e6981d1",
  2502 => x"cf029c74",
  2503 => x"4ba5c487",
  2504 => x"e2c37b74",
  2505 => x"f249bfd2",
  2506 => x"7b6e87c8",
  2507 => x"c4059c74",
  2508 => x"c24bc087",
  2509 => x"734bc187",
  2510 => x"87c9f249",
  2511 => x"c80266d4",
  2512 => x"eac04987",
  2513 => x"c24a7087",
  2514 => x"c24ac087",
  2515 => x"265aefdd",
  2516 => x"5887d7f1",
  2517 => x"1d141112",
  2518 => x"5a231c1b",
  2519 => x"f5949159",
  2520 => x"00f4ebf2",
  2521 => x"00000000",
  2522 => x"00000000",
  2523 => x"1e000000",
  2524 => x"c8ff4a71",
  2525 => x"a17249bf",
  2526 => x"1e4f2648",
  2527 => x"89bfc8ff",
  2528 => x"c0c0c0fe",
  2529 => x"01a9c0c0",
  2530 => x"4ac087c4",
  2531 => x"4ac187c2",
  2532 => x"4f264872",
  2533 => x"4ad4ff1e",
  2534 => x"c848d0ff",
  2535 => x"f0c378c5",
  2536 => x"c07a717a",
  2537 => x"7a7a7a7a",
  2538 => x"4f2678c4",
  2539 => x"4ad4ff1e",
  2540 => x"c848d0ff",
  2541 => x"7ac078c5",
  2542 => x"7ac0496a",
  2543 => x"7a7a7a7a",
  2544 => x"487178c4",
  2545 => x"5e0e4f26",
  2546 => x"0e5d5c5b",
  2547 => x"a6cc86e4",
  2548 => x"66ecc059",
  2549 => x"58a6dc48",
  2550 => x"e8c24d70",
  2551 => x"dae2c395",
  2552 => x"a5d8c285",
  2553 => x"48a6c47e",
  2554 => x"78a5dcc2",
  2555 => x"4cbf66c4",
  2556 => x"c294bf6e",
  2557 => x"946d85e0",
  2558 => x"c04b66c8",
  2559 => x"49c0c84a",
  2560 => x"87c1e3fd",
  2561 => x"c14866c8",
  2562 => x"c8789fc0",
  2563 => x"81c24966",
  2564 => x"799fbf6e",
  2565 => x"c64966c8",
  2566 => x"bf66c481",
  2567 => x"66c8799f",
  2568 => x"6d81cc49",
  2569 => x"66c8799f",
  2570 => x"d080d448",
  2571 => x"e3c258a6",
  2572 => x"66cc48ff",
  2573 => x"4aa1d449",
  2574 => x"aa714120",
  2575 => x"c887f905",
  2576 => x"eec04866",
  2577 => x"58a6d480",
  2578 => x"48d4e4c2",
  2579 => x"c84966d0",
  2580 => x"41204aa1",
  2581 => x"f905aa71",
  2582 => x"4866c887",
  2583 => x"d880f6c0",
  2584 => x"e4c258a6",
  2585 => x"66d448dd",
  2586 => x"a1e8c049",
  2587 => x"7141204a",
  2588 => x"87f905aa",
  2589 => x"c04a66d8",
  2590 => x"66d482f1",
  2591 => x"7281cb49",
  2592 => x"4966c851",
  2593 => x"c881dec1",
  2594 => x"799fd0c0",
  2595 => x"c14966c8",
  2596 => x"c0c881e2",
  2597 => x"66c8799f",
  2598 => x"81eac149",
  2599 => x"c8799fc1",
  2600 => x"ecc14966",
  2601 => x"9fbf6e81",
  2602 => x"4966c879",
  2603 => x"c481eec1",
  2604 => x"799fbf66",
  2605 => x"c14966c8",
  2606 => x"9f6d81f0",
  2607 => x"cf4b7479",
  2608 => x"739bffff",
  2609 => x"4966c84a",
  2610 => x"7281f2c1",
  2611 => x"4a74799f",
  2612 => x"ffcf2ad0",
  2613 => x"4c729aff",
  2614 => x"c14966c8",
  2615 => x"9f7481f4",
  2616 => x"66c87379",
  2617 => x"81f8c149",
  2618 => x"72799f73",
  2619 => x"c14966c8",
  2620 => x"9f7281fa",
  2621 => x"268ee479",
  2622 => x"264c264d",
  2623 => x"694f264b",
  2624 => x"6953544d",
  2625 => x"696e694d",
  2626 => x"7267484d",
  2627 => x"6c646661",
  2628 => x"00652069",
  2629 => x"3030312e",
  2630 => x"20202020",
  2631 => x"69446500",
  2632 => x"6653544d",
  2633 => x"20792069",
  2634 => x"20202020",
  2635 => x"20202020",
  2636 => x"20202020",
  2637 => x"20202020",
  2638 => x"20202020",
  2639 => x"20202020",
  2640 => x"20202020",
  2641 => x"731e0020",
  2642 => x"d44b711e",
  2643 => x"87d40266",
  2644 => x"d84966c8",
  2645 => x"c84a7331",
  2646 => x"49a17232",
  2647 => x"718166cc",
  2648 => x"87e3c048",
  2649 => x"c24966d0",
  2650 => x"e2c391e8",
  2651 => x"dcc281da",
  2652 => x"4a6a4aa1",
  2653 => x"66c89273",
  2654 => x"81e0c282",
  2655 => x"91724969",
  2656 => x"c18166cc",
  2657 => x"fd487189",
  2658 => x"711e87f1",
  2659 => x"49d4ff4a",
  2660 => x"c848d0ff",
  2661 => x"d0c278c5",
  2662 => x"7979c079",
  2663 => x"79797979",
  2664 => x"79727979",
  2665 => x"66c479c0",
  2666 => x"c879c079",
  2667 => x"79c07966",
  2668 => x"c07966cc",
  2669 => x"7966d079",
  2670 => x"66d479c0",
  2671 => x"2678c479",
  2672 => x"4a711e4f",
  2673 => x"9749a2c6",
  2674 => x"f0c34969",
  2675 => x"c01e7199",
  2676 => x"1ec11e1e",
  2677 => x"fe491ec0",
  2678 => x"d0c287f0",
  2679 => x"87f4f649",
  2680 => x"4f268eec",
  2681 => x"1e1ec01e",
  2682 => x"c11e1e1e",
  2683 => x"87dafe49",
  2684 => x"f649d0c2",
  2685 => x"8eec87de",
  2686 => x"711e4f26",
  2687 => x"48d0ff4a",
  2688 => x"ff78c5c8",
  2689 => x"e0c248d4",
  2690 => x"7878c078",
  2691 => x"c8787878",
  2692 => x"49721ec0",
  2693 => x"87dfdcfd",
  2694 => x"c448d0ff",
  2695 => x"4f262678",
  2696 => x"5c5b5e0e",
  2697 => x"86f80e5d",
  2698 => x"a2c24a71",
  2699 => x"7b97c14b",
  2700 => x"c14ca2c3",
  2701 => x"49a27c97",
  2702 => x"a2c451c0",
  2703 => x"7d97c04d",
  2704 => x"6e7ea2c5",
  2705 => x"c450c048",
  2706 => x"a2c648a6",
  2707 => x"4866c478",
  2708 => x"66d850c0",
  2709 => x"c6d1c31e",
  2710 => x"87eaf549",
  2711 => x"bf9766c8",
  2712 => x"66c81e49",
  2713 => x"1e49bf97",
  2714 => x"141e4915",
  2715 => x"49131e49",
  2716 => x"fc49c01e",
  2717 => x"49c887d4",
  2718 => x"c387d9f4",
  2719 => x"fd49c6d1",
  2720 => x"49d087f8",
  2721 => x"e087cdf4",
  2722 => x"87ebf98e",
  2723 => x"c64a711e",
  2724 => x"699749a2",
  2725 => x"a2c51e49",
  2726 => x"49699749",
  2727 => x"49a2c41e",
  2728 => x"1e496997",
  2729 => x"9749a2c3",
  2730 => x"c21e4969",
  2731 => x"699749a2",
  2732 => x"49c01e49",
  2733 => x"c287d3fb",
  2734 => x"d7f349d0",
  2735 => x"268eec87",
  2736 => x"1e731e4f",
  2737 => x"a2c24a71",
  2738 => x"d04b1149",
  2739 => x"c806abb7",
  2740 => x"49d1c287",
  2741 => x"d587fdf2",
  2742 => x"4966c887",
  2743 => x"c391e8c2",
  2744 => x"c281dae2",
  2745 => x"797381e4",
  2746 => x"f249d0c2",
  2747 => x"caf887e6",
  2748 => x"1e731e87",
  2749 => x"a3c64b71",
  2750 => x"49699749",
  2751 => x"49a3c51e",
  2752 => x"1e496997",
  2753 => x"9749a3c4",
  2754 => x"c31e4969",
  2755 => x"699749a3",
  2756 => x"a3c21e49",
  2757 => x"49699749",
  2758 => x"4aa3c11e",
  2759 => x"e9f94912",
  2760 => x"49d0c287",
  2761 => x"ec87edf1",
  2762 => x"87cff78e",
  2763 => x"5c5b5e0e",
  2764 => x"711e0e5d",
  2765 => x"c2496e7e",
  2766 => x"7997c181",
  2767 => x"83c34b6e",
  2768 => x"6e7b97c1",
  2769 => x"c082c14a",
  2770 => x"4c6e7a97",
  2771 => x"97c084c4",
  2772 => x"c54d6e7c",
  2773 => x"6e55c085",
  2774 => x"9785c64d",
  2775 => x"c01e4d6d",
  2776 => x"4c6c971e",
  2777 => x"4b6b971e",
  2778 => x"4969971e",
  2779 => x"f849121e",
  2780 => x"d0c287d8",
  2781 => x"87dcf049",
  2782 => x"faf58ee8",
  2783 => x"5b5e0e87",
  2784 => x"ff0e5d5c",
  2785 => x"4c7186dc",
  2786 => x"1149a4c3",
  2787 => x"4aa4c44d",
  2788 => x"9749a4c5",
  2789 => x"31c84969",
  2790 => x"484a6a97",
  2791 => x"a6d4b071",
  2792 => x"7ea4c658",
  2793 => x"49bf976e",
  2794 => x"d898cf48",
  2795 => x"487158a6",
  2796 => x"dc98c0c1",
  2797 => x"ec4858a6",
  2798 => x"78a4c280",
  2799 => x"bf9766c4",
  2800 => x"c3059b4b",
  2801 => x"4bc0c487",
  2802 => x"c01e66d8",
  2803 => x"751e66f8",
  2804 => x"66e0c01e",
  2805 => x"66e0c01e",
  2806 => x"87eaf549",
  2807 => x"497086d0",
  2808 => x"59a6e0c0",
  2809 => x"c5029b73",
  2810 => x"f8c087fb",
  2811 => x"87c50266",
  2812 => x"c55ba6d0",
  2813 => x"48a6cc87",
  2814 => x"66cc78c1",
  2815 => x"66f8c04c",
  2816 => x"c087de02",
  2817 => x"c24966f4",
  2818 => x"e2c391e8",
  2819 => x"e4c281da",
  2820 => x"48a6c881",
  2821 => x"66cc7869",
  2822 => x"b766c848",
  2823 => x"87c106a8",
  2824 => x"66fcc04c",
  2825 => x"c887d905",
  2826 => x"87e8ed49",
  2827 => x"7087fded",
  2828 => x"0599c449",
  2829 => x"f3ed87ca",
  2830 => x"c4497087",
  2831 => x"87f60299",
  2832 => x"88c14874",
  2833 => x"7058a6d0",
  2834 => x"029c744a",
  2835 => x"c187d4c1",
  2836 => x"c2c102ab",
  2837 => x"66f4c087",
  2838 => x"91e8c249",
  2839 => x"48dae2c3",
  2840 => x"a6cc8071",
  2841 => x"4966c858",
  2842 => x"6981e0c2",
  2843 => x"e4c005ad",
  2844 => x"d44dc187",
  2845 => x"80c14866",
  2846 => x"c858a6d8",
  2847 => x"dcc24966",
  2848 => x"05a86981",
  2849 => x"a6d487d1",
  2850 => x"d078c048",
  2851 => x"80c14866",
  2852 => x"c258a6d4",
  2853 => x"c185c187",
  2854 => x"c149728b",
  2855 => x"0599718a",
  2856 => x"d887ecfe",
  2857 => x"87d90266",
  2858 => x"66dc4974",
  2859 => x"c34a7181",
  2860 => x"4d729aff",
  2861 => x"b7c84a71",
  2862 => x"5aa6d42a",
  2863 => x"a629b7d8",
  2864 => x"bf976e59",
  2865 => x"99f0c349",
  2866 => x"71b166d4",
  2867 => x"4966d41e",
  2868 => x"7129b7c8",
  2869 => x"1e66d81e",
  2870 => x"66d41e75",
  2871 => x"1e49bf97",
  2872 => x"e5f249c0",
  2873 => x"c086d487",
  2874 => x"c10566fc",
  2875 => x"49d087f1",
  2876 => x"c087e1ea",
  2877 => x"c24966f4",
  2878 => x"e2c391e8",
  2879 => x"807148da",
  2880 => x"c858a6cc",
  2881 => x"81c84966",
  2882 => x"cdc10269",
  2883 => x"4966dc87",
  2884 => x"1e7131c9",
  2885 => x"fd4966cc",
  2886 => x"c487e5f8",
  2887 => x"a6e0c086",
  2888 => x"7866cc48",
  2889 => x"c0029c74",
  2890 => x"1ec087f5",
  2891 => x"fd4966cc",
  2892 => x"c187dbf2",
  2893 => x"4966d01e",
  2894 => x"87f1f0fd",
  2895 => x"66dc86c8",
  2896 => x"c080c148",
  2897 => x"c058a6e0",
  2898 => x"484966e0",
  2899 => x"e4c088c1",
  2900 => x"997158a6",
  2901 => x"87d2ff05",
  2902 => x"49c987c5",
  2903 => x"7387f5e8",
  2904 => x"c5fa059b",
  2905 => x"66fcc087",
  2906 => x"d087c502",
  2907 => x"87e4e849",
  2908 => x"ee8edcff",
  2909 => x"5e0e87c1",
  2910 => x"0e5d5c5b",
  2911 => x"4c7186e0",
  2912 => x"1149a4c3",
  2913 => x"58a6d448",
  2914 => x"c54aa4c4",
  2915 => x"699749a4",
  2916 => x"9731c849",
  2917 => x"71484a6a",
  2918 => x"58a6d8b0",
  2919 => x"6e7ea4c6",
  2920 => x"4d49bf97",
  2921 => x"48719dcf",
  2922 => x"dc98c0c1",
  2923 => x"ec4858a6",
  2924 => x"78a4c280",
  2925 => x"bf9766c4",
  2926 => x"1e66d84b",
  2927 => x"1e66f4c0",
  2928 => x"751e66d8",
  2929 => x"66e4c01e",
  2930 => x"87faed49",
  2931 => x"497086d0",
  2932 => x"59a6e0c0",
  2933 => x"c3059b73",
  2934 => x"4bc0c487",
  2935 => x"f3e649c4",
  2936 => x"4966dc87",
  2937 => x"1e7131c9",
  2938 => x"4966f4c0",
  2939 => x"c391e8c2",
  2940 => x"7148dae2",
  2941 => x"58a6d480",
  2942 => x"fd4966d0",
  2943 => x"c487c1f5",
  2944 => x"029b7386",
  2945 => x"c087dfc4",
  2946 => x"c40266f4",
  2947 => x"c24a7387",
  2948 => x"724ac187",
  2949 => x"66f4c04c",
  2950 => x"cc87d302",
  2951 => x"e4c24966",
  2952 => x"48a6c881",
  2953 => x"66c87869",
  2954 => x"c106aab7",
  2955 => x"9c744c87",
  2956 => x"87d5c202",
  2957 => x"7087f5e5",
  2958 => x"0599c849",
  2959 => x"ebe587ca",
  2960 => x"c8497087",
  2961 => x"87f60299",
  2962 => x"c848d0ff",
  2963 => x"d4ff78c5",
  2964 => x"78f0c248",
  2965 => x"787878c0",
  2966 => x"c0c87878",
  2967 => x"c6d1c31e",
  2968 => x"e8cbfd49",
  2969 => x"48d0ff87",
  2970 => x"d1c378c4",
  2971 => x"66d41ec6",
  2972 => x"dceefd49",
  2973 => x"d81ec187",
  2974 => x"ebfd4966",
  2975 => x"86cc87ef",
  2976 => x"c14866dc",
  2977 => x"a6e0c080",
  2978 => x"02abc158",
  2979 => x"cc87f3c0",
  2980 => x"e0c24966",
  2981 => x"4866d081",
  2982 => x"dd05a869",
  2983 => x"48a6d087",
  2984 => x"cc8578c1",
  2985 => x"dcc24966",
  2986 => x"05ad6981",
  2987 => x"4dc087d4",
  2988 => x"c14866d4",
  2989 => x"58a6d880",
  2990 => x"66d087c8",
  2991 => x"d480c148",
  2992 => x"8bc158a6",
  2993 => x"ebfd058c",
  2994 => x"0266d887",
  2995 => x"66dc87da",
  2996 => x"99ffc349",
  2997 => x"dc59a6d4",
  2998 => x"b7c84966",
  2999 => x"59a6d829",
  3000 => x"d84966dc",
  3001 => x"4d7129b7",
  3002 => x"49bf976e",
  3003 => x"7599f0c3",
  3004 => x"d81e71b1",
  3005 => x"b7c84966",
  3006 => x"dc1e7129",
  3007 => x"66dc1e66",
  3008 => x"9766d41e",
  3009 => x"c01e49bf",
  3010 => x"87fee949",
  3011 => x"9b7386d4",
  3012 => x"d087c702",
  3013 => x"87fce149",
  3014 => x"d0c287c6",
  3015 => x"87f4e149",
  3016 => x"fb059b73",
  3017 => x"8ee087e1",
  3018 => x"0e87cce7",
  3019 => x"5d5c5b5e",
  3020 => x"7186f80e",
  3021 => x"49a4c84c",
  3022 => x"2ac94a69",
  3023 => x"c3029a72",
  3024 => x"1e7287ca",
  3025 => x"4ad14972",
  3026 => x"87c6c6fd",
  3027 => x"99714a26",
  3028 => x"87c4c205",
  3029 => x"c0c0c4c1",
  3030 => x"fbc101aa",
  3031 => x"cc7ed187",
  3032 => x"01aac0f0",
  3033 => x"4dc487c5",
  3034 => x"7287ccc1",
  3035 => x"c649721e",
  3036 => x"ddc5fd4a",
  3037 => x"714a2687",
  3038 => x"87cc0599",
  3039 => x"aac0e0d9",
  3040 => x"c687c501",
  3041 => x"87efc04d",
  3042 => x"1e724bc5",
  3043 => x"4a734972",
  3044 => x"87fec4fd",
  3045 => x"99714a26",
  3046 => x"7387cb05",
  3047 => x"c0d0c449",
  3048 => x"06aa7191",
  3049 => x"abc587cf",
  3050 => x"c187c205",
  3051 => x"d083c183",
  3052 => x"d5ff04ab",
  3053 => x"724d7387",
  3054 => x"7549721e",
  3055 => x"d1c4fd4a",
  3056 => x"26497087",
  3057 => x"721e714a",
  3058 => x"fd4ad11e",
  3059 => x"2687c3c4",
  3060 => x"c849264a",
  3061 => x"87db58a6",
  3062 => x"d07effc0",
  3063 => x"c449724d",
  3064 => x"721e7129",
  3065 => x"4affc01e",
  3066 => x"87e6c3fd",
  3067 => x"49264a26",
  3068 => x"c258a6c8",
  3069 => x"c449a4d8",
  3070 => x"dcc27966",
  3071 => x"797549a4",
  3072 => x"49a4e0c2",
  3073 => x"e4c2796e",
  3074 => x"79c149a4",
  3075 => x"e6e38ef8",
  3076 => x"49c01e87",
  3077 => x"bfe2e2c3",
  3078 => x"c187c202",
  3079 => x"cae5c349",
  3080 => x"87c202bf",
  3081 => x"d0ffb1c2",
  3082 => x"78c5c848",
  3083 => x"c348d4ff",
  3084 => x"787178fa",
  3085 => x"c448d0ff",
  3086 => x"1e4f2678",
  3087 => x"4a711e73",
  3088 => x"4966cc1e",
  3089 => x"c391e8c2",
  3090 => x"714bdae2",
  3091 => x"fd497383",
  3092 => x"c487eee1",
  3093 => x"02987086",
  3094 => x"497387cb",
  3095 => x"87f3eafd",
  3096 => x"c6fb4973",
  3097 => x"87e9fe87",
  3098 => x"0e87d0e2",
  3099 => x"5d5c5b5e",
  3100 => x"ff86f40e",
  3101 => x"7087f5dc",
  3102 => x"0299c449",
  3103 => x"ff87ecc5",
  3104 => x"c5c848d0",
  3105 => x"48d4ff78",
  3106 => x"c078c0c2",
  3107 => x"78787878",
  3108 => x"d4ff4d78",
  3109 => x"7678c048",
  3110 => x"ff49a54a",
  3111 => x"7997bfd4",
  3112 => x"c048d4ff",
  3113 => x"c1516878",
  3114 => x"adb7c885",
  3115 => x"ff87e304",
  3116 => x"78c448d0",
  3117 => x"486697c6",
  3118 => x"7058a6cc",
  3119 => x"c49bd04b",
  3120 => x"49732bb7",
  3121 => x"c391e8c2",
  3122 => x"c881dae2",
  3123 => x"ca056981",
  3124 => x"49d1c287",
  3125 => x"87fcdaff",
  3126 => x"c787d0c4",
  3127 => x"494c6697",
  3128 => x"d099f0c3",
  3129 => x"87cc05a9",
  3130 => x"49721e73",
  3131 => x"c487d2e3",
  3132 => x"87f7c386",
  3133 => x"05acd0c2",
  3134 => x"497287c8",
  3135 => x"c387e5e3",
  3136 => x"ecc387e9",
  3137 => x"87ce05ac",
  3138 => x"1e731ec0",
  3139 => x"cfe44972",
  3140 => x"c386c887",
  3141 => x"d1c287d5",
  3142 => x"87cc05ac",
  3143 => x"49721e73",
  3144 => x"c487e9e5",
  3145 => x"87c3c386",
  3146 => x"05acc6c3",
  3147 => x"1e7387cc",
  3148 => x"cce64972",
  3149 => x"c286c487",
  3150 => x"e0c087f1",
  3151 => x"87cf05ac",
  3152 => x"731e1ec0",
  3153 => x"e849721e",
  3154 => x"86cc87f3",
  3155 => x"c387dcc2",
  3156 => x"d005acc4",
  3157 => x"c11ec087",
  3158 => x"721e731e",
  3159 => x"87dde849",
  3160 => x"c6c286cc",
  3161 => x"acf0c087",
  3162 => x"c087ce05",
  3163 => x"721e731e",
  3164 => x"87c2f049",
  3165 => x"f2c186c8",
  3166 => x"acc5c387",
  3167 => x"c187ce05",
  3168 => x"721e731e",
  3169 => x"87eeef49",
  3170 => x"dec186c8",
  3171 => x"05acc887",
  3172 => x"1e7387cc",
  3173 => x"d3e64972",
  3174 => x"c186c487",
  3175 => x"c0c187cd",
  3176 => x"87d005ac",
  3177 => x"1ec01ec1",
  3178 => x"49721e73",
  3179 => x"cc87cee7",
  3180 => x"87f7c086",
  3181 => x"cc059c74",
  3182 => x"721e7387",
  3183 => x"87f1e449",
  3184 => x"e6c086c4",
  3185 => x"1e66c887",
  3186 => x"496697c9",
  3187 => x"6697cc1e",
  3188 => x"97cf1e49",
  3189 => x"d21e4966",
  3190 => x"1e496697",
  3191 => x"deff49c4",
  3192 => x"86d487e8",
  3193 => x"ff49d1c2",
  3194 => x"f487e9d6",
  3195 => x"c6dcff8e",
  3196 => x"5b5e0e87",
  3197 => x"1e0e5d5c",
  3198 => x"d4ff7e71",
  3199 => x"c31e6e4b",
  3200 => x"fd49eae7",
  3201 => x"c487fada",
  3202 => x"9d4d7086",
  3203 => x"87c3c302",
  3204 => x"bff2e7c3",
  3205 => x"fd496e4c",
  3206 => x"ff87ddf6",
  3207 => x"c5c848d0",
  3208 => x"7bd6c178",
  3209 => x"7b154ac0",
  3210 => x"e0c082c1",
  3211 => x"f504aab7",
  3212 => x"48d0ff87",
  3213 => x"c5c878c4",
  3214 => x"7bd3c178",
  3215 => x"78c47bc1",
  3216 => x"c1029c74",
  3217 => x"d1c387fc",
  3218 => x"c0c87ec6",
  3219 => x"b7c08c4d",
  3220 => x"87c603ac",
  3221 => x"4da4c0c8",
  3222 => x"ddc34cc0",
  3223 => x"49bf97f7",
  3224 => x"d20299d0",
  3225 => x"c31ec087",
  3226 => x"fd49eae7",
  3227 => x"c487dfdd",
  3228 => x"4a497086",
  3229 => x"c387efc0",
  3230 => x"c31ec6d1",
  3231 => x"fd49eae7",
  3232 => x"c487cbdd",
  3233 => x"4a497086",
  3234 => x"c848d0ff",
  3235 => x"d4c178c5",
  3236 => x"bf976e7b",
  3237 => x"c1486e7b",
  3238 => x"c17e7080",
  3239 => x"f0ff058d",
  3240 => x"48d0ff87",
  3241 => x"9a7278c4",
  3242 => x"c087c505",
  3243 => x"87e5c048",
  3244 => x"e7c31ec1",
  3245 => x"dafd49ea",
  3246 => x"86c487f3",
  3247 => x"fe059c74",
  3248 => x"d0ff87c4",
  3249 => x"78c5c848",
  3250 => x"c07bd3c1",
  3251 => x"c178c47b",
  3252 => x"c087c248",
  3253 => x"4d262648",
  3254 => x"4b264c26",
  3255 => x"5e0e4f26",
  3256 => x"710e5c5b",
  3257 => x"0266cc4b",
  3258 => x"c04c87d8",
  3259 => x"d8028cf0",
  3260 => x"c14a7487",
  3261 => x"87d1028a",
  3262 => x"87cd028a",
  3263 => x"87c9028a",
  3264 => x"497387d0",
  3265 => x"c987eafb",
  3266 => x"731e7487",
  3267 => x"87ebf449",
  3268 => x"c3ff86c4",
  3269 => x"c31e0087",
  3270 => x"49bfe4cd",
  3271 => x"cdc3b9c1",
  3272 => x"d4ff59e8",
  3273 => x"78ffc348",
  3274 => x"c848d0ff",
  3275 => x"d4ff78e1",
  3276 => x"c478c148",
  3277 => x"ff787131",
  3278 => x"e0c048d0",
  3279 => x"1e4f2678",
  3280 => x"1ed8cdc3",
  3281 => x"49eae7c3",
  3282 => x"87f5d5fd",
  3283 => x"987086c4",
  3284 => x"ff87c302",
  3285 => x"4f2687c0",
  3286 => x"484b3531",
  3287 => x"2020205a",
  3288 => x"00474643",
  3289 => x"00000000",
  3290 => x"ede1c31e",
  3291 => x"b0c148bf",
  3292 => x"58f1e1c3",
  3293 => x"87d1e9fe",
  3294 => x"48d5ccc3",
  3295 => x"cfc350c2",
  3296 => x"f949bfd1",
  3297 => x"ccc387eb",
  3298 => x"50c148d5",
  3299 => x"bfcdcfc3",
  3300 => x"87ddf949",
  3301 => x"48d5ccc3",
  3302 => x"cfc350c3",
  3303 => x"f949bfd5",
  3304 => x"f0c087cf",
  3305 => x"d9cfc31e",
  3306 => x"f1fc49bf",
  3307 => x"1ef1c087",
  3308 => x"bfddcfc3",
  3309 => x"87e6fc49",
  3310 => x"bfede1c3",
  3311 => x"c398fe48",
  3312 => x"fe58f1e1",
  3313 => x"c087c2e8",
  3314 => x"268ef848",
  3315 => x"0033e14f",
  3316 => x"0033ed00",
  3317 => x"0033f900",
  3318 => x"00340500",
  3319 => x"00341100",
  3320 => x"58435000",
  3321 => x"20202054",
  3322 => x"4d4f5220",
  3323 => x"4e415400",
  3324 => x"20205944",
  3325 => x"4d4f5220",
  3326 => x"49545800",
  3327 => x"20204544",
  3328 => x"4d4f5220",
  3329 => x"58435000",
  3330 => x"20203154",
  3331 => x"44485620",
  3332 => x"58435000",
  3333 => x"20203254",
  3334 => x"44485620",
  3335 => x"44485600",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
